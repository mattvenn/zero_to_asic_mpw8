VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_simon_game
  CLASS BLOCK ;
  FOREIGN wrapped_simon_game ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 278.540 4.000 279.740 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.330 1.000 93.890 4.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.390 296.000 167.950 299.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.170 296.000 3.730 299.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 251.340 299.000 252.540 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.630 1.000 142.190 4.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.650 296.000 113.210 299.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 261.540 299.000 262.740 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 23.540 299.000 24.740 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.350 296.000 64.910 299.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.010 296.000 74.570 299.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.550 1.000 258.110 4.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 98.340 4.000 99.540 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 173.140 4.000 174.340 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 115.340 4.000 116.540 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 91.540 299.000 92.740 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.910 296.000 58.470 299.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.810 296.000 42.370 299.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.350 1.000 225.910 4.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.910 1.000 219.470 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 64.340 299.000 65.540 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.370 1.000 196.930 4.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.410 296.000 299.970 299.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.550 1.000 97.110 4.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 115.340 299.000 116.540 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 264.940 4.000 266.140 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.710 1.000 187.270 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 156.140 4.000 157.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.570 296.000 229.130 299.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.770 296.000 261.330 299.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 186.740 299.000 187.940 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.210 296.000 267.770 299.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 296.000 174.390 299.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 179.940 299.000 181.140 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 285.340 299.000 286.540 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 183.340 4.000 184.540 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 125.540 4.000 126.740 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 196.940 299.000 198.140 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.470 296.000 52.030 299.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.730 1.000 158.290 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 101.740 4.000 102.940 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 169.740 299.000 170.940 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 88.140 299.000 89.340 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 81.340 299.000 82.540 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 26.940 4.000 28.140 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.890 296.000 87.450 299.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 9.940 299.000 11.140 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.450 1.000 81.010 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.910 296.000 219.470 299.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.110 296.000 90.670 299.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.010 1.000 235.570 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 128.940 299.000 130.140 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.830 296.000 13.390 299.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 1.000 32.710 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.290 296.000 151.850 299.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.730 296.000 158.290 299.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.530 1.000 287.090 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 234.340 299.000 235.540 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.270 296.000 180.830 299.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.110 1.000 251.670 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 193.540 299.000 194.740 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.110 296.000 251.670 299.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.270 296.000 19.830 299.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.890 1.000 248.450 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 149.340 4.000 150.540 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.970 1.000 293.530 4.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 296.000 68.130 299.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 132.340 4.000 133.540 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 67.740 4.000 68.940 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 108.540 4.000 109.740 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.510 1.000 155.070 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 -0.260 299.000 0.940 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 196.940 4.000 198.140 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 105.140 299.000 106.340 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.450 296.000 81.010 299.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.710 1.000 26.270 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.350 1.000 64.910 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 278.540 299.000 279.740 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 162.940 299.000 164.140 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 16.740 4.000 17.940 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 43.940 4.000 45.140 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.450 1.000 242.010 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 237.740 299.000 238.940 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 247.940 4.000 249.140 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 156.140 299.000 157.340 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.090 296.000 280.650 299.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.090 1.000 280.650 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 142.540 4.000 143.740 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.810 296.000 203.370 299.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.670 296.000 245.230 299.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 244.540 4.000 245.740 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.150 1.000 193.710 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 132.340 299.000 133.540 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.170 1.000 164.730 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.130 296.000 222.690 299.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 33.740 4.000 34.940 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.010 296.000 235.570 299.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.990 1.000 103.550 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 6.540 299.000 7.740 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.810 1.000 42.370 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 40.540 4.000 41.740 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 84.740 4.000 85.940 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 285.340 4.000 286.540 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 40.540 299.000 41.740 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 244.540 299.000 245.740 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 227.540 299.000 228.740 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.550 296.000 97.110 299.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 268.340 299.000 269.540 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 261.540 4.000 262.740 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 173.140 299.000 174.340 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.630 296.000 142.190 299.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.750 296.000 290.310 299.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 122.140 4.000 123.340 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.870 1.000 116.430 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 91.540 4.000 92.740 ;
    END
  END io_out[9]
  PIN la1_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 47.340 299.000 48.540 ;
    END
  END la1_data_in[0]
  PIN la1_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.970 1.000 132.530 4.000 ;
    END
  END la1_data_in[10]
  PIN la1_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 33.740 299.000 34.940 ;
    END
  END la1_data_in[11]
  PIN la1_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 224.140 4.000 225.340 ;
    END
  END la1_data_in[12]
  PIN la1_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.810 1.000 203.370 4.000 ;
    END
  END la1_data_in[13]
  PIN la1_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 81.340 4.000 82.540 ;
    END
  END la1_data_in[14]
  PIN la1_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.990 296.000 103.550 299.000 ;
    END
  END la1_data_in[15]
  PIN la1_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.930 296.000 190.490 299.000 ;
    END
  END la1_data_in[16]
  PIN la1_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.850 296.000 145.410 299.000 ;
    END
  END la1_data_in[17]
  PIN la1_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.990 1.000 264.550 4.000 ;
    END
  END la1_data_in[18]
  PIN la1_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.210 296.000 106.770 299.000 ;
    END
  END la1_data_in[19]
  PIN la1_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.090 1.000 119.650 4.000 ;
    END
  END la1_data_in[1]
  PIN la1_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 220.740 4.000 221.940 ;
    END
  END la1_data_in[20]
  PIN la1_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.190 296.000 296.750 299.000 ;
    END
  END la1_data_in[21]
  PIN la1_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 50.740 299.000 51.940 ;
    END
  END la1_data_in[22]
  PIN la1_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 3.140 4.000 4.340 ;
    END
  END la1_data_in[23]
  PIN la1_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.890 1.000 87.450 4.000 ;
    END
  END la1_data_in[24]
  PIN la1_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 230.940 4.000 232.140 ;
    END
  END la1_data_in[25]
  PIN la1_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 16.740 299.000 17.940 ;
    END
  END la1_data_in[26]
  PIN la1_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 1.000 174.390 4.000 ;
    END
  END la1_data_in[27]
  PIN la1_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 203.740 4.000 204.940 ;
    END
  END la1_data_in[28]
  PIN la1_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.390 296.000 6.950 299.000 ;
    END
  END la1_data_in[29]
  PIN la1_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.790 1.000 71.350 4.000 ;
    END
  END la1_data_in[2]
  PIN la1_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.610 1.000 10.170 4.000 ;
    END
  END la1_data_in[30]
  PIN la1_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.790 1.000 232.350 4.000 ;
    END
  END la1_data_in[31]
  PIN la1_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 190.140 4.000 191.340 ;
    END
  END la1_data_in[3]
  PIN la1_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.550 296.000 258.110 299.000 ;
    END
  END la1_data_in[4]
  PIN la1_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 145.940 299.000 147.140 ;
    END
  END la1_data_in[5]
  PIN la1_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.090 296.000 119.650 299.000 ;
    END
  END la1_data_in[6]
  PIN la1_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 139.140 4.000 140.340 ;
    END
  END la1_data_in[7]
  PIN la1_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.530 296.000 126.090 299.000 ;
    END
  END la1_data_in[8]
  PIN la1_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 207.140 4.000 208.340 ;
    END
  END la1_data_in[9]
  PIN la1_data_out[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.250 1.000 48.810 4.000 ;
    END
  END la1_data_out[0]
  PIN la1_data_out[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 71.140 299.000 72.340 ;
    END
  END la1_data_out[10]
  PIN la1_data_out[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.190 1.000 135.750 4.000 ;
    END
  END la1_data_out[11]
  PIN la1_data_out[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 275.140 299.000 276.340 ;
    END
  END la1_data_out[12]
  PIN la1_data_out[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.930 296.000 29.490 299.000 ;
    END
  END la1_data_out[13]
  PIN la1_data_out[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.170 296.000 164.730 299.000 ;
    END
  END la1_data_out[14]
  PIN la1_data_out[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 9.940 4.000 11.140 ;
    END
  END la1_data_out[15]
  PIN la1_data_out[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 98.340 299.000 99.540 ;
    END
  END la1_data_out[16]
  PIN la1_data_out[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 213.940 299.000 215.140 ;
    END
  END la1_data_out[17]
  PIN la1_data_out[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.370 296.000 35.930 299.000 ;
    END
  END la1_data_out[18]
  PIN la1_data_out[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 152.740 299.000 153.940 ;
    END
  END la1_data_out[19]
  PIN la1_data_out[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 271.740 4.000 272.940 ;
    END
  END la1_data_out[1]
  PIN la1_data_out[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 60.940 4.000 62.140 ;
    END
  END la1_data_out[20]
  PIN la1_data_out[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 254.740 299.000 255.940 ;
    END
  END la1_data_out[21]
  PIN la1_data_out[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.490 296.000 184.050 299.000 ;
    END
  END la1_data_out[22]
  PIN la1_data_out[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.230 1.000 77.790 4.000 ;
    END
  END la1_data_out[23]
  PIN la1_data_out[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 111.940 299.000 113.140 ;
    END
  END la1_data_out[24]
  PIN la1_data_out[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 20.140 4.000 21.340 ;
    END
  END la1_data_out[25]
  PIN la1_data_out[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 30.340 299.000 31.540 ;
    END
  END la1_data_out[26]
  PIN la1_data_out[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 288.740 4.000 289.940 ;
    END
  END la1_data_out[27]
  PIN la1_data_out[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.430 1.000 270.990 4.000 ;
    END
  END la1_data_out[28]
  PIN la1_data_out[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.590 1.000 39.150 4.000 ;
    END
  END la1_data_out[29]
  PIN la1_data_out[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.530 1.000 126.090 4.000 ;
    END
  END la1_data_out[2]
  PIN la1_data_out[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 74.540 299.000 75.740 ;
    END
  END la1_data_out[30]
  PIN la1_data_out[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 292.140 299.000 293.340 ;
    END
  END la1_data_out[31]
  PIN la1_data_out[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 57.540 4.000 58.740 ;
    END
  END la1_data_out[3]
  PIN la1_data_out[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.650 1.000 274.210 4.000 ;
    END
  END la1_data_out[4]
  PIN la1_data_out[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.270 1.000 19.830 4.000 ;
    END
  END la1_data_out[5]
  PIN la1_data_out[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 122.140 299.000 123.340 ;
    END
  END la1_data_out[6]
  PIN la1_data_out[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.170 1.000 3.730 4.000 ;
    END
  END la1_data_out[7]
  PIN la1_data_out[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 220.740 299.000 221.940 ;
    END
  END la1_data_out[8]
  PIN la1_data_out[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.310 296.000 283.870 299.000 ;
    END
  END la1_data_out[9]
  PIN la1_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.190 1.000 296.750 4.000 ;
    END
  END la1_oenb[0]
  PIN la1_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.650 296.000 274.210 299.000 ;
    END
  END la1_oenb[10]
  PIN la1_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 166.340 4.000 167.540 ;
    END
  END la1_oenb[11]
  PIN la1_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 179.940 4.000 181.140 ;
    END
  END la1_oenb[12]
  PIN la1_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.270 1.000 180.830 4.000 ;
    END
  END la1_oenb[13]
  PIN la1_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 1.000 0.510 4.000 ;
    END
  END la1_oenb[14]
  PIN la1_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.470 1.000 213.030 4.000 ;
    END
  END la1_oenb[15]
  PIN la1_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 213.940 4.000 215.140 ;
    END
  END la1_oenb[16]
  PIN la1_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.710 296.000 26.270 299.000 ;
    END
  END la1_oenb[17]
  PIN la1_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.190 296.000 135.750 299.000 ;
    END
  END la1_oenb[18]
  PIN la1_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 162.940 4.000 164.140 ;
    END
  END la1_oenb[19]
  PIN la1_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.690 1.000 55.250 4.000 ;
    END
  END la1_oenb[1]
  PIN la1_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.050 1.000 16.610 4.000 ;
    END
  END la1_oenb[20]
  PIN la1_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.370 296.000 196.930 299.000 ;
    END
  END la1_oenb[21]
  PIN la1_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.750 296.000 129.310 299.000 ;
    END
  END la1_oenb[22]
  PIN la1_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.070 1.000 148.630 4.000 ;
    END
  END la1_oenb[23]
  PIN la1_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.450 296.000 242.010 299.000 ;
    END
  END la1_oenb[24]
  PIN la1_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 57.540 299.000 58.740 ;
    END
  END la1_oenb[25]
  PIN la1_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 237.740 4.000 238.940 ;
    END
  END la1_oenb[26]
  PIN la1_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 210.540 299.000 211.740 ;
    END
  END la1_oenb[27]
  PIN la1_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.910 1.000 58.470 4.000 ;
    END
  END la1_oenb[28]
  PIN la1_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.430 1.000 109.990 4.000 ;
    END
  END la1_oenb[29]
  PIN la1_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 50.740 4.000 51.940 ;
    END
  END la1_oenb[2]
  PIN la1_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 203.740 299.000 204.940 ;
    END
  END la1_oenb[30]
  PIN la1_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.610 1.000 171.170 4.000 ;
    END
  END la1_oenb[31]
  PIN la1_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.470 296.000 213.030 299.000 ;
    END
  END la1_oenb[3]
  PIN la1_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.030 296.000 206.590 299.000 ;
    END
  END la1_oenb[4]
  PIN la1_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 295.540 4.000 296.740 ;
    END
  END la1_oenb[5]
  PIN la1_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.250 296.000 48.810 299.000 ;
    END
  END la1_oenb[6]
  PIN la1_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.250 1.000 209.810 4.000 ;
    END
  END la1_oenb[7]
  PIN la1_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 74.540 4.000 75.740 ;
    END
  END la1_oenb[8]
  PIN la1_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 254.740 4.000 255.940 ;
    END
  END la1_oenb[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 139.140 299.000 140.340 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 294.400 288.405 ;
      LAYER met1 ;
        RECT 3.290 10.640 294.400 288.560 ;
      LAYER met2 ;
        RECT 4.010 295.720 6.110 296.000 ;
        RECT 7.230 295.720 12.550 296.000 ;
        RECT 13.670 295.720 18.990 296.000 ;
        RECT 20.110 295.720 25.430 296.000 ;
        RECT 26.550 295.720 28.650 296.000 ;
        RECT 29.770 295.720 35.090 296.000 ;
        RECT 36.210 295.720 41.530 296.000 ;
        RECT 42.650 295.720 47.970 296.000 ;
        RECT 49.090 295.720 51.190 296.000 ;
        RECT 52.310 295.720 57.630 296.000 ;
        RECT 58.750 295.720 64.070 296.000 ;
        RECT 65.190 295.720 67.290 296.000 ;
        RECT 68.410 295.720 73.730 296.000 ;
        RECT 74.850 295.720 80.170 296.000 ;
        RECT 81.290 295.720 86.610 296.000 ;
        RECT 87.730 295.720 89.830 296.000 ;
        RECT 90.950 295.720 96.270 296.000 ;
        RECT 97.390 295.720 102.710 296.000 ;
        RECT 103.830 295.720 105.930 296.000 ;
        RECT 107.050 295.720 112.370 296.000 ;
        RECT 113.490 295.720 118.810 296.000 ;
        RECT 119.930 295.720 125.250 296.000 ;
        RECT 126.370 295.720 128.470 296.000 ;
        RECT 129.590 295.720 134.910 296.000 ;
        RECT 136.030 295.720 141.350 296.000 ;
        RECT 142.470 295.720 144.570 296.000 ;
        RECT 145.690 295.720 151.010 296.000 ;
        RECT 152.130 295.720 157.450 296.000 ;
        RECT 158.570 295.720 163.890 296.000 ;
        RECT 165.010 295.720 167.110 296.000 ;
        RECT 168.230 295.720 173.550 296.000 ;
        RECT 174.670 295.720 179.990 296.000 ;
        RECT 181.110 295.720 183.210 296.000 ;
        RECT 184.330 295.720 189.650 296.000 ;
        RECT 190.770 295.720 196.090 296.000 ;
        RECT 197.210 295.720 202.530 296.000 ;
        RECT 203.650 295.720 205.750 296.000 ;
        RECT 206.870 295.720 212.190 296.000 ;
        RECT 213.310 295.720 218.630 296.000 ;
        RECT 219.750 295.720 221.850 296.000 ;
        RECT 222.970 295.720 228.290 296.000 ;
        RECT 229.410 295.720 234.730 296.000 ;
        RECT 235.850 295.720 241.170 296.000 ;
        RECT 242.290 295.720 244.390 296.000 ;
        RECT 245.510 295.720 250.830 296.000 ;
        RECT 251.950 295.720 257.270 296.000 ;
        RECT 258.390 295.720 260.490 296.000 ;
        RECT 261.610 295.720 266.930 296.000 ;
        RECT 268.050 295.720 273.370 296.000 ;
        RECT 274.490 295.720 279.810 296.000 ;
        RECT 280.930 295.720 283.030 296.000 ;
        RECT 284.150 295.720 289.470 296.000 ;
        RECT 290.590 295.720 293.380 296.000 ;
        RECT 3.320 4.280 293.380 295.720 ;
        RECT 4.010 0.720 9.330 4.280 ;
        RECT 10.450 0.720 15.770 4.280 ;
        RECT 16.890 0.720 18.990 4.280 ;
        RECT 20.110 0.720 25.430 4.280 ;
        RECT 26.550 0.720 31.870 4.280 ;
        RECT 32.990 0.720 38.310 4.280 ;
        RECT 39.430 0.720 41.530 4.280 ;
        RECT 42.650 0.720 47.970 4.280 ;
        RECT 49.090 0.720 54.410 4.280 ;
        RECT 55.530 0.720 57.630 4.280 ;
        RECT 58.750 0.720 64.070 4.280 ;
        RECT 65.190 0.720 70.510 4.280 ;
        RECT 71.630 0.720 76.950 4.280 ;
        RECT 78.070 0.720 80.170 4.280 ;
        RECT 81.290 0.720 86.610 4.280 ;
        RECT 87.730 0.720 93.050 4.280 ;
        RECT 94.170 0.720 96.270 4.280 ;
        RECT 97.390 0.720 102.710 4.280 ;
        RECT 103.830 0.720 109.150 4.280 ;
        RECT 110.270 0.720 115.590 4.280 ;
        RECT 116.710 0.720 118.810 4.280 ;
        RECT 119.930 0.720 125.250 4.280 ;
        RECT 126.370 0.720 131.690 4.280 ;
        RECT 132.810 0.720 134.910 4.280 ;
        RECT 136.030 0.720 141.350 4.280 ;
        RECT 142.470 0.720 147.790 4.280 ;
        RECT 148.910 0.720 154.230 4.280 ;
        RECT 155.350 0.720 157.450 4.280 ;
        RECT 158.570 0.720 163.890 4.280 ;
        RECT 165.010 0.720 170.330 4.280 ;
        RECT 171.450 0.720 173.550 4.280 ;
        RECT 174.670 0.720 179.990 4.280 ;
        RECT 181.110 0.720 186.430 4.280 ;
        RECT 187.550 0.720 192.870 4.280 ;
        RECT 193.990 0.720 196.090 4.280 ;
        RECT 197.210 0.720 202.530 4.280 ;
        RECT 203.650 0.720 208.970 4.280 ;
        RECT 210.090 0.720 212.190 4.280 ;
        RECT 213.310 0.720 218.630 4.280 ;
        RECT 219.750 0.720 225.070 4.280 ;
        RECT 226.190 0.720 231.510 4.280 ;
        RECT 232.630 0.720 234.730 4.280 ;
        RECT 235.850 0.720 241.170 4.280 ;
        RECT 242.290 0.720 247.610 4.280 ;
        RECT 248.730 0.720 250.830 4.280 ;
        RECT 251.950 0.720 257.270 4.280 ;
        RECT 258.390 0.720 263.710 4.280 ;
        RECT 264.830 0.720 270.150 4.280 ;
        RECT 271.270 0.720 273.370 4.280 ;
        RECT 274.490 0.720 279.810 4.280 ;
        RECT 280.930 0.720 286.250 4.280 ;
        RECT 287.370 0.720 292.690 4.280 ;
        RECT 3.320 0.155 293.380 0.720 ;
      LAYER met3 ;
        RECT 4.000 291.740 295.600 292.905 ;
        RECT 4.000 290.340 296.000 291.740 ;
        RECT 4.400 288.340 296.000 290.340 ;
        RECT 4.000 286.940 296.000 288.340 ;
        RECT 4.400 284.940 295.600 286.940 ;
        RECT 4.000 280.140 296.000 284.940 ;
        RECT 4.400 278.140 295.600 280.140 ;
        RECT 4.000 276.740 296.000 278.140 ;
        RECT 4.000 274.740 295.600 276.740 ;
        RECT 4.000 273.340 296.000 274.740 ;
        RECT 4.400 271.340 296.000 273.340 ;
        RECT 4.000 269.940 296.000 271.340 ;
        RECT 4.000 267.940 295.600 269.940 ;
        RECT 4.000 266.540 296.000 267.940 ;
        RECT 4.400 264.540 296.000 266.540 ;
        RECT 4.000 263.140 296.000 264.540 ;
        RECT 4.400 261.140 295.600 263.140 ;
        RECT 4.000 256.340 296.000 261.140 ;
        RECT 4.400 254.340 295.600 256.340 ;
        RECT 4.000 252.940 296.000 254.340 ;
        RECT 4.000 250.940 295.600 252.940 ;
        RECT 4.000 249.540 296.000 250.940 ;
        RECT 4.400 247.540 296.000 249.540 ;
        RECT 4.000 246.140 296.000 247.540 ;
        RECT 4.400 244.140 295.600 246.140 ;
        RECT 4.000 239.340 296.000 244.140 ;
        RECT 4.400 237.340 295.600 239.340 ;
        RECT 4.000 235.940 296.000 237.340 ;
        RECT 4.000 233.940 295.600 235.940 ;
        RECT 4.000 232.540 296.000 233.940 ;
        RECT 4.400 230.540 296.000 232.540 ;
        RECT 4.000 229.140 296.000 230.540 ;
        RECT 4.000 227.140 295.600 229.140 ;
        RECT 4.000 225.740 296.000 227.140 ;
        RECT 4.400 223.740 296.000 225.740 ;
        RECT 4.000 222.340 296.000 223.740 ;
        RECT 4.400 220.340 295.600 222.340 ;
        RECT 4.000 215.540 296.000 220.340 ;
        RECT 4.400 213.540 295.600 215.540 ;
        RECT 4.000 212.140 296.000 213.540 ;
        RECT 4.000 210.140 295.600 212.140 ;
        RECT 4.000 208.740 296.000 210.140 ;
        RECT 4.400 206.740 296.000 208.740 ;
        RECT 4.000 205.340 296.000 206.740 ;
        RECT 4.400 203.340 295.600 205.340 ;
        RECT 4.000 198.540 296.000 203.340 ;
        RECT 4.400 196.540 295.600 198.540 ;
        RECT 4.000 195.140 296.000 196.540 ;
        RECT 4.000 193.140 295.600 195.140 ;
        RECT 4.000 191.740 296.000 193.140 ;
        RECT 4.400 189.740 296.000 191.740 ;
        RECT 4.000 188.340 296.000 189.740 ;
        RECT 4.000 186.340 295.600 188.340 ;
        RECT 4.000 184.940 296.000 186.340 ;
        RECT 4.400 182.940 296.000 184.940 ;
        RECT 4.000 181.540 296.000 182.940 ;
        RECT 4.400 179.540 295.600 181.540 ;
        RECT 4.000 174.740 296.000 179.540 ;
        RECT 4.400 172.740 295.600 174.740 ;
        RECT 4.000 171.340 296.000 172.740 ;
        RECT 4.000 169.340 295.600 171.340 ;
        RECT 4.000 167.940 296.000 169.340 ;
        RECT 4.400 165.940 296.000 167.940 ;
        RECT 4.000 164.540 296.000 165.940 ;
        RECT 4.400 162.540 295.600 164.540 ;
        RECT 4.000 157.740 296.000 162.540 ;
        RECT 4.400 155.740 295.600 157.740 ;
        RECT 4.000 154.340 296.000 155.740 ;
        RECT 4.000 152.340 295.600 154.340 ;
        RECT 4.000 150.940 296.000 152.340 ;
        RECT 4.400 148.940 296.000 150.940 ;
        RECT 4.000 147.540 296.000 148.940 ;
        RECT 4.000 145.540 295.600 147.540 ;
        RECT 4.000 144.140 296.000 145.540 ;
        RECT 4.400 142.140 296.000 144.140 ;
        RECT 4.000 140.740 296.000 142.140 ;
        RECT 4.400 138.740 295.600 140.740 ;
        RECT 4.000 133.940 296.000 138.740 ;
        RECT 4.400 131.940 295.600 133.940 ;
        RECT 4.000 130.540 296.000 131.940 ;
        RECT 4.000 128.540 295.600 130.540 ;
        RECT 4.000 127.140 296.000 128.540 ;
        RECT 4.400 125.140 296.000 127.140 ;
        RECT 4.000 123.740 296.000 125.140 ;
        RECT 4.400 121.740 295.600 123.740 ;
        RECT 4.000 116.940 296.000 121.740 ;
        RECT 4.400 114.940 295.600 116.940 ;
        RECT 4.000 113.540 296.000 114.940 ;
        RECT 4.000 111.540 295.600 113.540 ;
        RECT 4.000 110.140 296.000 111.540 ;
        RECT 4.400 108.140 296.000 110.140 ;
        RECT 4.000 106.740 296.000 108.140 ;
        RECT 4.000 104.740 295.600 106.740 ;
        RECT 4.000 103.340 296.000 104.740 ;
        RECT 4.400 101.340 296.000 103.340 ;
        RECT 4.000 99.940 296.000 101.340 ;
        RECT 4.400 97.940 295.600 99.940 ;
        RECT 4.000 93.140 296.000 97.940 ;
        RECT 4.400 91.140 295.600 93.140 ;
        RECT 4.000 89.740 296.000 91.140 ;
        RECT 4.000 87.740 295.600 89.740 ;
        RECT 4.000 86.340 296.000 87.740 ;
        RECT 4.400 84.340 296.000 86.340 ;
        RECT 4.000 82.940 296.000 84.340 ;
        RECT 4.400 80.940 295.600 82.940 ;
        RECT 4.000 76.140 296.000 80.940 ;
        RECT 4.400 74.140 295.600 76.140 ;
        RECT 4.000 72.740 296.000 74.140 ;
        RECT 4.000 70.740 295.600 72.740 ;
        RECT 4.000 69.340 296.000 70.740 ;
        RECT 4.400 67.340 296.000 69.340 ;
        RECT 4.000 65.940 296.000 67.340 ;
        RECT 4.000 63.940 295.600 65.940 ;
        RECT 4.000 62.540 296.000 63.940 ;
        RECT 4.400 60.540 296.000 62.540 ;
        RECT 4.000 59.140 296.000 60.540 ;
        RECT 4.400 57.140 295.600 59.140 ;
        RECT 4.000 52.340 296.000 57.140 ;
        RECT 4.400 50.340 295.600 52.340 ;
        RECT 4.000 48.940 296.000 50.340 ;
        RECT 4.000 46.940 295.600 48.940 ;
        RECT 4.000 45.540 296.000 46.940 ;
        RECT 4.400 43.540 296.000 45.540 ;
        RECT 4.000 42.140 296.000 43.540 ;
        RECT 4.400 40.140 295.600 42.140 ;
        RECT 4.000 35.340 296.000 40.140 ;
        RECT 4.400 33.340 295.600 35.340 ;
        RECT 4.000 31.940 296.000 33.340 ;
        RECT 4.000 29.940 295.600 31.940 ;
        RECT 4.000 28.540 296.000 29.940 ;
        RECT 4.400 26.540 296.000 28.540 ;
        RECT 4.000 25.140 296.000 26.540 ;
        RECT 4.000 23.140 295.600 25.140 ;
        RECT 4.000 21.740 296.000 23.140 ;
        RECT 4.400 19.740 296.000 21.740 ;
        RECT 4.000 18.340 296.000 19.740 ;
        RECT 4.400 16.340 295.600 18.340 ;
        RECT 4.000 11.540 296.000 16.340 ;
        RECT 4.400 9.540 295.600 11.540 ;
        RECT 4.000 8.140 296.000 9.540 ;
        RECT 4.000 6.140 295.600 8.140 ;
        RECT 4.000 4.740 296.000 6.140 ;
        RECT 4.400 2.740 296.000 4.740 ;
        RECT 4.000 1.340 296.000 2.740 ;
        RECT 4.000 0.175 295.600 1.340 ;
      LAYER met4 ;
        RECT 85.855 46.415 97.440 267.065 ;
        RECT 99.840 46.415 174.240 267.065 ;
        RECT 176.640 46.415 235.225 267.065 ;
  END
END wrapped_simon_game
END LIBRARY

