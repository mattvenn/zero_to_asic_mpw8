magic
tech sky130A
magscale 1 2
timestamp 1672435764
<< metal1 >>
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 188338 700476 188344 700528
rect 188396 700516 188402 700528
rect 267642 700516 267648 700528
rect 188396 700488 267648 700516
rect 188396 700476 188402 700488
rect 267642 700476 267648 700488
rect 267700 700476 267706 700528
rect 40494 700408 40500 700460
rect 40552 700448 40558 700460
rect 78674 700448 78680 700460
rect 40552 700420 78680 700448
rect 40552 700408 40558 700420
rect 78674 700408 78680 700420
rect 78732 700408 78738 700460
rect 89162 700408 89168 700460
rect 89220 700448 89226 700460
rect 122834 700448 122840 700460
rect 89220 700420 122840 700448
rect 89220 700408 89226 700420
rect 122834 700408 122840 700420
rect 122892 700408 122898 700460
rect 184198 700408 184204 700460
rect 184256 700448 184262 700460
rect 364978 700448 364984 700460
rect 184256 700420 364984 700448
rect 184256 700408 184262 700420
rect 364978 700408 364984 700420
rect 365036 700408 365042 700460
rect 73062 700340 73068 700392
rect 73120 700380 73126 700392
rect 137830 700380 137836 700392
rect 73120 700352 137836 700380
rect 73120 700340 73126 700352
rect 137830 700340 137836 700352
rect 137888 700340 137894 700392
rect 182818 700340 182824 700392
rect 182876 700380 182882 700392
rect 429838 700380 429844 700392
rect 182876 700352 429844 700380
rect 182876 700340 182882 700352
rect 429838 700340 429844 700352
rect 429896 700340 429902 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 94498 700312 94504 700324
rect 8168 700284 94504 700312
rect 8168 700272 8174 700284
rect 94498 700272 94504 700284
rect 94556 700272 94562 700324
rect 105446 700272 105452 700324
rect 105504 700312 105510 700324
rect 120718 700312 120724 700324
rect 105504 700284 120724 700312
rect 105504 700272 105510 700284
rect 120718 700272 120724 700284
rect 120776 700272 120782 700324
rect 186958 700272 186964 700324
rect 187016 700312 187022 700324
rect 527174 700312 527180 700324
rect 187016 700284 527180 700312
rect 187016 700272 187022 700284
rect 527174 700272 527180 700284
rect 527232 700272 527238 700324
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 25498 699700 25504 699712
rect 24360 699672 25504 699700
rect 24360 699660 24366 699672
rect 25498 699660 25504 699672
rect 25556 699660 25562 699712
rect 66162 699660 66168 699712
rect 66220 699700 66226 699712
rect 72970 699700 72976 699712
rect 66220 699672 72976 699700
rect 66220 699660 66226 699672
rect 72970 699660 72976 699672
rect 73028 699660 73034 699712
rect 396718 699660 396724 699712
rect 396776 699700 396782 699712
rect 397454 699700 397460 699712
rect 396776 699672 397460 699700
rect 396776 699660 396782 699672
rect 397454 699660 397460 699672
rect 397512 699660 397518 699712
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 75914 683176 75920 683188
rect 3476 683148 75920 683176
rect 3476 683136 3482 683148
rect 75914 683136 75920 683148
rect 75972 683136 75978 683188
rect 233878 683136 233884 683188
rect 233936 683176 233942 683188
rect 579614 683176 579620 683188
rect 233936 683148 579620 683176
rect 233936 683136 233942 683148
rect 579614 683136 579620 683148
rect 579672 683136 579678 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 55858 670732 55864 670744
rect 3568 670704 55864 670732
rect 3568 670692 3574 670704
rect 55858 670692 55864 670704
rect 55916 670692 55922 670744
rect 192478 670692 192484 670744
rect 192536 670732 192542 670744
rect 580166 670732 580172 670744
rect 192536 670704 580172 670732
rect 192536 670692 192542 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 95878 656928 95884 656940
rect 3476 656900 95884 656928
rect 3476 656888 3482 656900
rect 95878 656888 95884 656900
rect 95936 656888 95942 656940
rect 249058 643084 249064 643136
rect 249116 643124 249122 643136
rect 580166 643124 580172 643136
rect 249116 643096 580172 643124
rect 249116 643084 249122 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 54478 632108 54484 632120
rect 3476 632080 54484 632108
rect 3476 632068 3482 632080
rect 54478 632068 54484 632080
rect 54536 632068 54542 632120
rect 239398 630640 239404 630692
rect 239456 630680 239462 630692
rect 579982 630680 579988 630692
rect 239456 630652 579988 630680
rect 239456 630640 239462 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 106274 618304 106280 618316
rect 3200 618276 106280 618304
rect 3200 618264 3206 618276
rect 106274 618264 106280 618276
rect 106332 618264 106338 618316
rect 235258 616836 235264 616888
rect 235316 616876 235322 616888
rect 580166 616876 580172 616888
rect 235316 616848 580172 616876
rect 235316 616836 235322 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 62758 605860 62764 605872
rect 3292 605832 62764 605860
rect 3292 605820 3298 605832
rect 62758 605820 62764 605832
rect 62816 605820 62822 605872
rect 242158 590656 242164 590708
rect 242216 590696 242222 590708
rect 580166 590696 580172 590708
rect 242216 590668 580172 590696
rect 242216 590656 242222 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 65518 579680 65524 579692
rect 3384 579652 65524 579680
rect 3384 579640 3390 579652
rect 65518 579640 65524 579652
rect 65576 579640 65582 579692
rect 169662 576852 169668 576904
rect 169720 576892 169726 576904
rect 580166 576892 580172 576904
rect 169720 576864 580172 576892
rect 169720 576852 169726 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 11698 565876 11704 565888
rect 3476 565848 11704 565876
rect 3476 565836 3482 565848
rect 11698 565836 11704 565848
rect 11756 565836 11762 565888
rect 233970 563048 233976 563100
rect 234028 563088 234034 563100
rect 580166 563088 580172 563100
rect 234028 563060 580172 563088
rect 234028 563048 234034 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 121454 553432 121460 553444
rect 3476 553404 121460 553432
rect 3476 553392 3482 553404
rect 121454 553392 121460 553404
rect 121512 553392 121518 553444
rect 278038 536800 278044 536852
rect 278096 536840 278102 536852
rect 579890 536840 579896 536852
rect 278096 536812 579896 536840
rect 278096 536800 278102 536812
rect 579890 536800 579896 536812
rect 579948 536800 579954 536852
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 120810 527184 120816 527196
rect 3476 527156 120816 527184
rect 3476 527144 3482 527156
rect 120810 527144 120816 527156
rect 120868 527144 120874 527196
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 107654 514808 107660 514820
rect 3476 514780 107660 514808
rect 3476 514768 3482 514780
rect 107654 514768 107660 514780
rect 107712 514768 107718 514820
rect 173158 510620 173164 510672
rect 173216 510660 173222 510672
rect 580166 510660 580172 510672
rect 173216 510632 580172 510660
rect 173216 510620 173222 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 99374 501004 99380 501016
rect 3108 500976 99380 501004
rect 3108 500964 3114 500976
rect 99374 500964 99380 500976
rect 99432 500964 99438 501016
rect 169570 484372 169576 484424
rect 169628 484412 169634 484424
rect 580166 484412 580172 484424
rect 169628 484384 580172 484412
rect 169628 484372 169634 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 2774 474784 2780 474836
rect 2832 474824 2838 474836
rect 4798 474824 4804 474836
rect 2832 474796 4804 474824
rect 2832 474784 2838 474796
rect 4798 474784 4804 474796
rect 4856 474784 4862 474836
rect 289078 470568 289084 470620
rect 289136 470608 289142 470620
rect 580166 470608 580172 470620
rect 289136 470580 580172 470608
rect 289136 470568 289142 470580
rect 580166 470568 580172 470580
rect 580224 470568 580230 470620
rect 3234 462340 3240 462392
rect 3292 462380 3298 462392
rect 18598 462380 18604 462392
rect 3292 462352 18604 462380
rect 3292 462340 3298 462352
rect 18598 462340 18604 462352
rect 18656 462340 18662 462392
rect 203518 456764 203524 456816
rect 203576 456804 203582 456816
rect 580166 456804 580172 456816
rect 203576 456776 580172 456804
rect 203576 456764 203582 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 61378 448576 61384 448588
rect 3200 448548 61384 448576
rect 3200 448536 3206 448548
rect 61378 448536 61384 448548
rect 61436 448536 61442 448588
rect 3418 422288 3424 422340
rect 3476 422328 3482 422340
rect 119338 422328 119344 422340
rect 3476 422300 119344 422328
rect 3476 422288 3482 422300
rect 119338 422288 119344 422300
rect 119396 422288 119402 422340
rect 169846 418140 169852 418192
rect 169904 418180 169910 418192
rect 580166 418180 580172 418192
rect 169904 418152 580172 418180
rect 169904 418140 169910 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 180058 404336 180064 404388
rect 180116 404376 180122 404388
rect 580166 404376 580172 404388
rect 180116 404348 580172 404376
rect 180116 404336 180122 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3510 397468 3516 397520
rect 3568 397508 3574 397520
rect 10318 397508 10324 397520
rect 3568 397480 10324 397508
rect 3568 397468 3574 397480
rect 10318 397468 10324 397480
rect 10376 397468 10382 397520
rect 238018 378156 238024 378208
rect 238076 378196 238082 378208
rect 580166 378196 580172 378208
rect 238076 378168 580172 378196
rect 238076 378156 238082 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 244918 364352 244924 364404
rect 244976 364392 244982 364404
rect 579798 364392 579804 364404
rect 244976 364364 579804 364392
rect 244976 364352 244982 364364
rect 579798 364352 579804 364364
rect 579856 364352 579862 364404
rect 234062 351908 234068 351960
rect 234120 351948 234126 351960
rect 580166 351948 580172 351960
rect 234120 351920 580172 351948
rect 234120 351908 234126 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 71774 345080 71780 345092
rect 3384 345052 71780 345080
rect 3384 345040 3390 345052
rect 71774 345040 71780 345052
rect 71832 345040 71838 345092
rect 195238 324300 195244 324352
rect 195296 324340 195302 324352
rect 579614 324340 579620 324352
rect 195296 324312 579620 324340
rect 195296 324300 195302 324312
rect 579614 324300 579620 324312
rect 579672 324300 579678 324352
rect 3326 318792 3332 318844
rect 3384 318832 3390 318844
rect 15838 318832 15844 318844
rect 3384 318804 15844 318832
rect 3384 318792 3390 318804
rect 15838 318792 15844 318804
rect 15896 318792 15902 318844
rect 169938 311856 169944 311908
rect 169996 311896 170002 311908
rect 580166 311896 580172 311908
rect 169996 311868 580172 311896
rect 169996 311856 170002 311868
rect 580166 311856 580172 311868
rect 580224 311856 580230 311908
rect 169018 298120 169024 298172
rect 169076 298160 169082 298172
rect 580166 298160 580172 298172
rect 169076 298132 580172 298160
rect 169076 298120 169082 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 3326 292544 3332 292596
rect 3384 292584 3390 292596
rect 58618 292584 58624 292596
rect 3384 292556 58624 292584
rect 3384 292544 3390 292556
rect 58618 292544 58624 292556
rect 58676 292544 58682 292596
rect 3418 266364 3424 266416
rect 3476 266404 3482 266416
rect 7558 266404 7564 266416
rect 3476 266376 7564 266404
rect 3476 266364 3482 266376
rect 7558 266364 7564 266376
rect 7616 266364 7622 266416
rect 123662 265616 123668 265668
rect 123720 265656 123726 265668
rect 201494 265656 201500 265668
rect 123720 265628 201500 265656
rect 123720 265616 123726 265628
rect 201494 265616 201500 265628
rect 201552 265616 201558 265668
rect 3602 260108 3608 260160
rect 3660 260148 3666 260160
rect 120166 260148 120172 260160
rect 3660 260120 120172 260148
rect 3660 260108 3666 260120
rect 120166 260108 120172 260120
rect 120224 260108 120230 260160
rect 3326 258680 3332 258732
rect 3384 258720 3390 258732
rect 120350 258720 120356 258732
rect 3384 258692 120356 258720
rect 3384 258680 3390 258692
rect 120350 258680 120356 258692
rect 120408 258680 120414 258732
rect 228358 258068 228364 258120
rect 228416 258108 228422 258120
rect 579982 258108 579988 258120
rect 228416 258080 579988 258108
rect 228416 258068 228422 258080
rect 579982 258068 579988 258080
rect 580040 258068 580046 258120
rect 25498 257320 25504 257372
rect 25556 257360 25562 257372
rect 121914 257360 121920 257372
rect 25556 257332 121920 257360
rect 25556 257320 25562 257332
rect 121914 257320 121920 257332
rect 121972 257320 121978 257372
rect 167730 257320 167736 257372
rect 167788 257360 167794 257372
rect 542354 257360 542360 257372
rect 167788 257332 542360 257360
rect 167788 257320 167794 257332
rect 542354 257320 542360 257332
rect 542412 257320 542418 257372
rect 10318 255960 10324 256012
rect 10376 256000 10382 256012
rect 121730 256000 121736 256012
rect 10376 255972 121736 256000
rect 10376 255960 10382 255972
rect 121730 255960 121736 255972
rect 121788 255960 121794 256012
rect 170030 255960 170036 256012
rect 170088 256000 170094 256012
rect 234614 256000 234620 256012
rect 170088 255972 234620 256000
rect 170088 255960 170094 255972
rect 234614 255960 234620 255972
rect 234672 255960 234678 256012
rect 65886 254736 65892 254788
rect 65944 254776 65950 254788
rect 170030 254776 170036 254788
rect 65944 254748 170036 254776
rect 65944 254736 65950 254748
rect 170030 254736 170036 254748
rect 170088 254736 170094 254788
rect 104158 254668 104164 254720
rect 104216 254708 104222 254720
rect 155218 254708 155224 254720
rect 104216 254680 155224 254708
rect 104216 254668 104222 254680
rect 155218 254668 155224 254680
rect 155276 254668 155282 254720
rect 91278 254600 91284 254652
rect 91336 254640 91342 254652
rect 91336 254612 142154 254640
rect 91336 254600 91342 254612
rect 68738 254532 68744 254584
rect 68796 254572 68802 254584
rect 126330 254572 126336 254584
rect 68796 254544 126336 254572
rect 68796 254532 68802 254544
rect 126330 254532 126336 254544
rect 126388 254532 126394 254584
rect 142126 254572 142154 254612
rect 142890 254572 142896 254584
rect 142126 254544 142896 254572
rect 142890 254532 142896 254544
rect 142948 254572 142954 254584
rect 194594 254572 194600 254584
rect 142948 254544 194600 254572
rect 142948 254532 142954 254544
rect 194594 254532 194600 254544
rect 194652 254532 194658 254584
rect 91922 254464 91928 254516
rect 91980 254504 91986 254516
rect 151078 254504 151084 254516
rect 91980 254476 151084 254504
rect 91980 254464 91986 254476
rect 151078 254464 151084 254476
rect 151136 254504 151142 254516
rect 195974 254504 195980 254516
rect 151136 254476 195980 254504
rect 151136 254464 151142 254476
rect 195974 254464 195980 254476
rect 196032 254464 196038 254516
rect 67542 254396 67548 254448
rect 67600 254436 67606 254448
rect 153194 254436 153200 254448
rect 67600 254408 153200 254436
rect 67600 254396 67606 254408
rect 153194 254396 153200 254408
rect 153252 254436 153258 254448
rect 153838 254436 153844 254448
rect 153252 254408 153844 254436
rect 153252 254396 153258 254408
rect 153838 254396 153844 254408
rect 153896 254396 153902 254448
rect 69290 254328 69296 254380
rect 69348 254368 69354 254380
rect 167270 254368 167276 254380
rect 69348 254340 167276 254368
rect 69348 254328 69354 254340
rect 167270 254328 167276 254340
rect 167328 254328 167334 254380
rect 69014 254260 69020 254312
rect 69072 254300 69078 254312
rect 167178 254300 167184 254312
rect 69072 254272 167184 254300
rect 69072 254260 69078 254272
rect 167178 254260 167184 254272
rect 167236 254260 167242 254312
rect 69382 254192 69388 254244
rect 69440 254232 69446 254244
rect 167638 254232 167644 254244
rect 69440 254204 167644 254232
rect 69440 254192 69446 254204
rect 167638 254192 167644 254204
rect 167696 254192 167702 254244
rect 67450 254124 67456 254176
rect 67508 254164 67514 254176
rect 167730 254164 167736 254176
rect 67508 254136 167736 254164
rect 67508 254124 67514 254136
rect 167730 254124 167736 254136
rect 167788 254124 167794 254176
rect 73890 254056 73896 254108
rect 73948 254096 73954 254108
rect 173986 254096 173992 254108
rect 73948 254068 173992 254096
rect 73948 254056 73954 254068
rect 173986 254056 173992 254068
rect 174044 254056 174050 254108
rect 77754 253988 77760 254040
rect 77812 254028 77818 254040
rect 179414 254028 179420 254040
rect 77812 254000 179420 254028
rect 77812 253988 77818 254000
rect 179414 253988 179420 254000
rect 179472 253988 179478 254040
rect 3142 253920 3148 253972
rect 3200 253960 3206 253972
rect 10318 253960 10324 253972
rect 3200 253932 10324 253960
rect 3200 253920 3206 253932
rect 10318 253920 10324 253932
rect 10376 253920 10382 253972
rect 114462 253920 114468 253972
rect 114520 253960 114526 253972
rect 126974 253960 126980 253972
rect 114520 253932 126980 253960
rect 114520 253920 114526 253932
rect 126974 253920 126980 253932
rect 127032 253920 127038 253972
rect 155218 253920 155224 253972
rect 155276 253960 155282 253972
rect 211154 253960 211160 253972
rect 155276 253932 211160 253960
rect 155276 253920 155282 253932
rect 211154 253920 211160 253932
rect 211212 253920 211218 253972
rect 80974 253512 80980 253564
rect 81032 253552 81038 253564
rect 183646 253552 183652 253564
rect 81032 253524 183652 253552
rect 81032 253512 81038 253524
rect 183646 253512 183652 253524
rect 183704 253512 183710 253564
rect 68462 253444 68468 253496
rect 68520 253484 68526 253496
rect 124858 253484 124864 253496
rect 68520 253456 124864 253484
rect 68520 253444 68526 253456
rect 124858 253444 124864 253456
rect 124916 253444 124922 253496
rect 99006 253376 99012 253428
rect 99064 253416 99070 253428
rect 204898 253416 204904 253428
rect 99064 253388 204904 253416
rect 99064 253376 99070 253388
rect 204898 253376 204904 253388
rect 204956 253376 204962 253428
rect 93210 253240 93216 253292
rect 93268 253280 93274 253292
rect 126238 253280 126244 253292
rect 93268 253252 126244 253280
rect 93268 253240 93274 253252
rect 126238 253240 126244 253252
rect 126296 253280 126302 253292
rect 126882 253280 126888 253292
rect 126296 253252 126888 253280
rect 126296 253240 126302 253252
rect 126882 253240 126888 253252
rect 126940 253240 126946 253292
rect 85482 253172 85488 253224
rect 85540 253212 85546 253224
rect 133322 253212 133328 253224
rect 85540 253184 133328 253212
rect 85540 253172 85546 253184
rect 133322 253172 133328 253184
rect 133380 253172 133386 253224
rect 68738 253104 68744 253156
rect 68796 253144 68802 253156
rect 120902 253144 120908 253156
rect 68796 253116 120908 253144
rect 68796 253104 68802 253116
rect 120902 253104 120908 253116
rect 120960 253104 120966 253156
rect 93854 253036 93860 253088
rect 93912 253076 93918 253088
rect 148318 253076 148324 253088
rect 93912 253048 148324 253076
rect 93912 253036 93918 253048
rect 148318 253036 148324 253048
rect 148376 253076 148382 253088
rect 198734 253076 198740 253088
rect 148376 253048 198740 253076
rect 148376 253036 148382 253048
rect 198734 253036 198740 253048
rect 198792 253036 198798 253088
rect 68278 252968 68284 253020
rect 68336 253008 68342 253020
rect 124030 253008 124036 253020
rect 68336 252980 124036 253008
rect 68336 252968 68342 252980
rect 124030 252968 124036 252980
rect 124088 252968 124094 253020
rect 126882 252968 126888 253020
rect 126940 253008 126946 253020
rect 181438 253008 181444 253020
rect 126940 252980 181444 253008
rect 126940 252968 126946 252980
rect 181438 252968 181444 252980
rect 181496 252968 181502 253020
rect 90634 252900 90640 252952
rect 90692 252940 90698 252952
rect 164142 252940 164148 252952
rect 90692 252912 164148 252940
rect 90692 252900 90698 252912
rect 164142 252900 164148 252912
rect 164200 252940 164206 252952
rect 194686 252940 194692 252952
rect 164200 252912 194692 252940
rect 164200 252900 164206 252912
rect 194686 252900 194692 252912
rect 194744 252900 194750 252952
rect 111886 252832 111892 252884
rect 111944 252872 111950 252884
rect 142798 252872 142804 252884
rect 111944 252844 142804 252872
rect 111944 252832 111950 252844
rect 142798 252832 142804 252844
rect 142856 252872 142862 252884
rect 219434 252872 219440 252884
rect 142856 252844 219440 252872
rect 142856 252832 142862 252844
rect 219434 252832 219440 252844
rect 219492 252832 219498 252884
rect 89346 252764 89352 252816
rect 89404 252804 89410 252816
rect 165522 252804 165528 252816
rect 89404 252776 165528 252804
rect 89404 252764 89410 252776
rect 165522 252764 165528 252776
rect 165580 252804 165586 252816
rect 193214 252804 193220 252816
rect 165580 252776 193220 252804
rect 165580 252764 165586 252776
rect 193214 252764 193220 252776
rect 193272 252764 193278 252816
rect 69474 252696 69480 252748
rect 69532 252736 69538 252748
rect 167822 252736 167828 252748
rect 69532 252708 167828 252736
rect 69532 252696 69538 252708
rect 167822 252696 167828 252708
rect 167880 252696 167886 252748
rect 112530 252628 112536 252680
rect 112588 252668 112594 252680
rect 120994 252668 121000 252680
rect 112588 252640 121000 252668
rect 112588 252628 112594 252640
rect 120994 252628 121000 252640
rect 121052 252628 121058 252680
rect 103514 252560 103520 252612
rect 103572 252600 103578 252612
rect 119982 252600 119988 252612
rect 103572 252572 119988 252600
rect 103572 252560 103578 252572
rect 119982 252560 119988 252572
rect 120040 252560 120046 252612
rect 109954 252220 109960 252272
rect 110012 252260 110018 252272
rect 118050 252260 118056 252272
rect 110012 252232 118056 252260
rect 110012 252220 110018 252232
rect 118050 252220 118056 252232
rect 118108 252220 118114 252272
rect 105446 252152 105452 252204
rect 105504 252192 105510 252204
rect 118786 252192 118792 252204
rect 105504 252164 118792 252192
rect 105504 252152 105510 252164
rect 118786 252152 118792 252164
rect 118844 252152 118850 252204
rect 80330 252084 80336 252136
rect 80388 252124 80394 252136
rect 112162 252124 112168 252136
rect 80388 252096 112168 252124
rect 80388 252084 80394 252096
rect 112162 252084 112168 252096
rect 112220 252084 112226 252136
rect 113174 252084 113180 252136
rect 113232 252124 113238 252136
rect 124214 252124 124220 252136
rect 113232 252096 124220 252124
rect 113232 252084 113238 252096
rect 124214 252084 124220 252096
rect 124272 252084 124278 252136
rect 69198 252016 69204 252068
rect 69256 252056 69262 252068
rect 71774 252056 71780 252068
rect 69256 252028 71780 252056
rect 69256 252016 69262 252028
rect 71774 252016 71780 252028
rect 71832 252056 71838 252068
rect 72602 252056 72608 252068
rect 71832 252028 72608 252056
rect 71832 252016 71838 252028
rect 72602 252016 72608 252028
rect 72660 252056 72666 252068
rect 121362 252056 121368 252068
rect 72660 252028 121368 252056
rect 72660 252016 72666 252028
rect 121362 252016 121368 252028
rect 121420 252016 121426 252068
rect 102226 251948 102232 252000
rect 102284 251988 102290 252000
rect 157978 251988 157984 252000
rect 102284 251960 157984 251988
rect 102284 251948 102290 251960
rect 157978 251948 157984 251960
rect 158036 251948 158042 252000
rect 71314 251880 71320 251932
rect 71372 251920 71378 251932
rect 122098 251920 122104 251932
rect 71372 251892 122104 251920
rect 71372 251880 71378 251892
rect 122098 251880 122104 251892
rect 122156 251880 122162 251932
rect 75822 251812 75828 251864
rect 75880 251852 75886 251864
rect 130378 251852 130384 251864
rect 75880 251824 130384 251852
rect 75880 251812 75886 251824
rect 130378 251812 130384 251824
rect 130436 251812 130442 251864
rect 108022 251744 108028 251796
rect 108080 251784 108086 251796
rect 124306 251784 124312 251796
rect 108080 251756 124312 251784
rect 108080 251744 108086 251756
rect 124306 251744 124312 251756
rect 124364 251744 124370 251796
rect 101582 251676 101588 251728
rect 101640 251716 101646 251728
rect 125134 251716 125140 251728
rect 101640 251688 125140 251716
rect 101640 251676 101646 251688
rect 125134 251676 125140 251688
rect 125192 251676 125198 251728
rect 66070 251608 66076 251660
rect 66128 251648 66134 251660
rect 75914 251648 75920 251660
rect 66128 251620 75920 251648
rect 66128 251608 66134 251620
rect 75914 251608 75920 251620
rect 75972 251648 75978 251660
rect 76466 251648 76472 251660
rect 75972 251620 76472 251648
rect 75972 251608 75978 251620
rect 76466 251608 76472 251620
rect 76524 251648 76530 251660
rect 95142 251648 95148 251660
rect 76524 251620 95148 251648
rect 76524 251608 76530 251620
rect 95142 251608 95148 251620
rect 95200 251608 95206 251660
rect 97074 251608 97080 251660
rect 97132 251648 97138 251660
rect 127802 251648 127808 251660
rect 97132 251620 127808 251648
rect 97132 251608 97138 251620
rect 127802 251608 127808 251620
rect 127860 251608 127866 251660
rect 62022 251540 62028 251592
rect 62080 251580 62086 251592
rect 85482 251580 85488 251592
rect 62080 251552 85488 251580
rect 62080 251540 62086 251552
rect 85482 251540 85488 251552
rect 85540 251540 85546 251592
rect 86770 251540 86776 251592
rect 86828 251580 86834 251592
rect 124122 251580 124128 251592
rect 86828 251552 124128 251580
rect 86828 251540 86834 251552
rect 124122 251540 124128 251552
rect 124180 251540 124186 251592
rect 63402 251472 63408 251524
rect 63460 251512 63466 251524
rect 74534 251512 74540 251524
rect 63460 251484 74540 251512
rect 63460 251472 63466 251484
rect 74534 251472 74540 251484
rect 74592 251512 74598 251524
rect 122190 251512 122196 251524
rect 74592 251484 122196 251512
rect 74592 251472 74598 251484
rect 122190 251472 122196 251484
rect 122248 251472 122254 251524
rect 117038 251404 117044 251456
rect 117096 251444 117102 251456
rect 126698 251444 126704 251456
rect 117096 251416 126704 251444
rect 117096 251404 117102 251416
rect 126698 251404 126704 251416
rect 126756 251404 126762 251456
rect 61746 251336 61752 251388
rect 61804 251376 61810 251388
rect 80974 251376 80980 251388
rect 61804 251348 80980 251376
rect 61804 251336 61810 251348
rect 80974 251336 80980 251348
rect 81032 251336 81038 251388
rect 110598 251336 110604 251388
rect 110656 251376 110662 251388
rect 121270 251376 121276 251388
rect 110656 251348 121276 251376
rect 110656 251336 110662 251348
rect 121270 251336 121276 251348
rect 121328 251336 121334 251388
rect 157978 251336 157984 251388
rect 158036 251376 158042 251388
rect 177298 251376 177304 251388
rect 158036 251348 177304 251376
rect 158036 251336 158042 251348
rect 177298 251336 177304 251348
rect 177356 251336 177362 251388
rect 97718 251268 97724 251320
rect 97776 251308 97782 251320
rect 103422 251308 103428 251320
rect 97776 251280 103428 251308
rect 97776 251268 97782 251280
rect 103422 251268 103428 251280
rect 103480 251268 103486 251320
rect 118326 251268 118332 251320
rect 118384 251308 118390 251320
rect 144178 251308 144184 251320
rect 118384 251280 144184 251308
rect 118384 251268 118390 251280
rect 144178 251268 144184 251280
rect 144236 251308 144242 251320
rect 211062 251308 211068 251320
rect 144236 251280 211068 251308
rect 144236 251268 144242 251280
rect 211062 251268 211068 251280
rect 211120 251268 211126 251320
rect 61930 251200 61936 251252
rect 61988 251240 61994 251252
rect 75822 251240 75828 251252
rect 61988 251212 75828 251240
rect 61988 251200 61994 251212
rect 75822 251200 75828 251212
rect 75880 251200 75886 251252
rect 100294 251200 100300 251252
rect 100352 251240 100358 251252
rect 117222 251240 117228 251252
rect 100352 251212 117228 251240
rect 100352 251200 100358 251212
rect 117222 251200 117228 251212
rect 117280 251200 117286 251252
rect 118970 251200 118976 251252
rect 119028 251240 119034 251252
rect 126606 251240 126612 251252
rect 119028 251212 126612 251240
rect 119028 251200 119034 251212
rect 126606 251200 126612 251212
rect 126664 251200 126670 251252
rect 131114 251200 131120 251252
rect 131172 251240 131178 251252
rect 131850 251240 131856 251252
rect 131172 251212 131856 251240
rect 131172 251200 131178 251212
rect 131850 251200 131856 251212
rect 131908 251240 131914 251252
rect 222838 251240 222844 251252
rect 131908 251212 222844 251240
rect 131908 251200 131914 251212
rect 222838 251200 222844 251212
rect 222896 251200 222902 251252
rect 107654 251132 107660 251184
rect 107712 251172 107718 251184
rect 108666 251172 108672 251184
rect 107712 251144 108672 251172
rect 107712 251132 107718 251144
rect 108666 251132 108672 251144
rect 108724 251132 108730 251184
rect 203058 251132 203064 251184
rect 203116 251172 203122 251184
rect 203518 251172 203524 251184
rect 203116 251144 203524 251172
rect 203116 251132 203122 251144
rect 203518 251132 203524 251144
rect 203576 251132 203582 251184
rect 211062 251132 211068 251184
rect 211120 251172 211126 251184
rect 227714 251172 227720 251184
rect 211120 251144 227720 251172
rect 211120 251132 211126 251144
rect 227714 251132 227720 251144
rect 227772 251172 227778 251184
rect 228358 251172 228364 251184
rect 227772 251144 228364 251172
rect 227772 251132 227778 251144
rect 228358 251132 228364 251144
rect 228416 251132 228422 251184
rect 117958 250724 117964 250776
rect 118016 250764 118022 250776
rect 125042 250764 125048 250776
rect 118016 250736 125048 250764
rect 118016 250724 118022 250736
rect 125042 250724 125048 250736
rect 125100 250724 125106 250776
rect 68186 250656 68192 250708
rect 68244 250696 68250 250708
rect 123846 250696 123852 250708
rect 68244 250668 123852 250696
rect 68244 250656 68250 250668
rect 123846 250656 123852 250668
rect 123904 250656 123910 250708
rect 108666 250588 108672 250640
rect 108724 250628 108730 250640
rect 134518 250628 134524 250640
rect 108724 250600 134524 250628
rect 108724 250588 108730 250600
rect 134518 250588 134524 250600
rect 134576 250588 134582 250640
rect 95878 250520 95884 250572
rect 95936 250560 95942 250572
rect 95936 250532 103514 250560
rect 95936 250520 95942 250532
rect 103486 250492 103514 250532
rect 117222 250520 117228 250572
rect 117280 250560 117286 250572
rect 129734 250560 129740 250572
rect 117280 250532 129740 250560
rect 117280 250520 117286 250532
rect 129734 250520 129740 250532
rect 129792 250520 129798 250572
rect 130470 250492 130476 250504
rect 103486 250464 130476 250492
rect 130470 250452 130476 250464
rect 130528 250452 130534 250504
rect 82906 250384 82912 250436
rect 82964 250424 82970 250436
rect 121086 250424 121092 250436
rect 82964 250396 121092 250424
rect 82964 250384 82970 250396
rect 121086 250384 121092 250396
rect 121144 250384 121150 250436
rect 68002 250316 68008 250368
rect 68060 250356 68066 250368
rect 123938 250356 123944 250368
rect 68060 250328 123944 250356
rect 68060 250316 68066 250328
rect 123938 250316 123944 250328
rect 123996 250316 124002 250368
rect 68646 250248 68652 250300
rect 68704 250288 68710 250300
rect 124950 250288 124956 250300
rect 68704 250260 124956 250288
rect 68704 250248 68710 250260
rect 124950 250248 124956 250260
rect 125008 250248 125014 250300
rect 68830 250180 68836 250232
rect 68888 250220 68894 250232
rect 117958 250220 117964 250232
rect 68888 250192 117964 250220
rect 68888 250180 68894 250192
rect 117958 250180 117964 250192
rect 118016 250180 118022 250232
rect 127710 250152 127716 250164
rect 84166 250124 127716 250152
rect 67910 250044 67916 250096
rect 67968 250084 67974 250096
rect 84166 250084 84194 250124
rect 127710 250112 127716 250124
rect 127768 250112 127774 250164
rect 146938 250152 146944 250164
rect 142126 250124 146944 250152
rect 67968 250056 84194 250084
rect 67968 250044 67974 250056
rect 87414 250044 87420 250096
rect 87472 250084 87478 250096
rect 142126 250084 142154 250124
rect 146938 250112 146944 250124
rect 146996 250152 147002 250164
rect 190454 250152 190460 250164
rect 146996 250124 190460 250152
rect 146996 250112 147002 250124
rect 190454 250112 190460 250124
rect 190512 250112 190518 250164
rect 87472 250056 142154 250084
rect 87472 250044 87478 250056
rect 152458 250044 152464 250096
rect 152516 250084 152522 250096
rect 203058 250084 203064 250096
rect 152516 250056 203064 250084
rect 152516 250044 152522 250056
rect 203058 250044 203064 250056
rect 203116 250044 203122 250096
rect 63310 249976 63316 250028
rect 63368 250016 63374 250028
rect 82906 250016 82912 250028
rect 63368 249988 82912 250016
rect 63368 249976 63374 249988
rect 82906 249976 82912 249988
rect 82964 249976 82970 250028
rect 99650 249976 99656 250028
rect 99708 250016 99714 250028
rect 121178 250016 121184 250028
rect 99708 249988 121184 250016
rect 99708 249976 99714 249988
rect 121178 249976 121184 249988
rect 121236 249976 121242 250028
rect 129734 249976 129740 250028
rect 129792 250016 129798 250028
rect 130562 250016 130568 250028
rect 129792 249988 130568 250016
rect 129792 249976 129798 249988
rect 130562 249976 130568 249988
rect 130620 250016 130626 250028
rect 205726 250016 205732 250028
rect 130620 249988 205732 250016
rect 130620 249976 130626 249988
rect 205726 249976 205732 249988
rect 205784 249976 205790 250028
rect 68370 249908 68376 249960
rect 68428 249948 68434 249960
rect 123478 249948 123484 249960
rect 68428 249920 123484 249948
rect 68428 249908 68434 249920
rect 123478 249908 123484 249920
rect 123536 249908 123542 249960
rect 130470 249908 130476 249960
rect 130528 249948 130534 249960
rect 201494 249948 201500 249960
rect 130528 249920 201500 249948
rect 130528 249908 130534 249920
rect 201494 249908 201500 249920
rect 201552 249908 201558 249960
rect 106734 249840 106740 249892
rect 106792 249880 106798 249892
rect 140038 249880 140044 249892
rect 106792 249852 140044 249880
rect 106792 249840 106798 249852
rect 140038 249840 140044 249852
rect 140096 249880 140102 249892
rect 210418 249880 210424 249892
rect 140096 249852 210424 249880
rect 140096 249840 140102 249852
rect 210418 249840 210424 249852
rect 210476 249840 210482 249892
rect 64782 249772 64788 249824
rect 64840 249812 64846 249824
rect 78674 249812 78680 249824
rect 64840 249784 78680 249812
rect 64840 249772 64846 249784
rect 78674 249772 78680 249784
rect 78732 249812 78738 249824
rect 79226 249812 79232 249824
rect 78732 249784 79232 249812
rect 78732 249772 78738 249784
rect 79226 249772 79232 249784
rect 79284 249812 79290 249824
rect 119798 249812 119804 249824
rect 79284 249784 119804 249812
rect 79284 249772 79290 249784
rect 119798 249772 119804 249784
rect 119856 249772 119862 249824
rect 134518 249772 134524 249824
rect 134576 249812 134582 249824
rect 215938 249812 215944 249824
rect 134576 249784 215944 249812
rect 134576 249772 134582 249784
rect 215938 249772 215944 249784
rect 215996 249772 216002 249824
rect 118694 249704 118700 249756
rect 118752 249744 118758 249756
rect 187694 249744 187700 249756
rect 118752 249716 187700 249744
rect 118752 249704 118758 249716
rect 187694 249704 187700 249716
rect 187752 249744 187758 249756
rect 188338 249744 188344 249756
rect 187752 249716 188344 249744
rect 187752 249704 187758 249716
rect 188338 249704 188344 249716
rect 188396 249704 188402 249756
rect 119154 249636 119160 249688
rect 119212 249676 119218 249688
rect 119430 249676 119436 249688
rect 119212 249648 119436 249676
rect 119212 249636 119218 249648
rect 119430 249636 119436 249648
rect 119488 249636 119494 249688
rect 115474 249500 115480 249552
rect 115532 249540 115538 249552
rect 119154 249540 119160 249552
rect 115532 249512 119160 249540
rect 115532 249500 115538 249512
rect 119154 249500 119160 249512
rect 119212 249500 119218 249552
rect 118050 249432 118056 249484
rect 118108 249432 118114 249484
rect 118786 249432 118792 249484
rect 118844 249472 118850 249484
rect 118844 249444 122834 249472
rect 118844 249432 118850 249444
rect 67082 249092 67088 249144
rect 67140 249132 67146 249144
rect 67542 249132 67548 249144
rect 67140 249104 67548 249132
rect 67140 249092 67146 249104
rect 67542 249092 67548 249104
rect 67600 249092 67606 249144
rect 118068 249064 118096 249432
rect 119706 249092 119712 249144
rect 119764 249132 119770 249144
rect 121546 249132 121552 249144
rect 119764 249104 121552 249132
rect 119764 249092 119770 249104
rect 121546 249092 121552 249104
rect 121604 249092 121610 249144
rect 122806 249132 122834 249444
rect 156598 249132 156604 249144
rect 122806 249104 156604 249132
rect 156598 249092 156604 249104
rect 156656 249092 156662 249144
rect 159358 249064 159364 249076
rect 118068 249036 159364 249064
rect 159358 249024 159364 249036
rect 159416 249024 159422 249076
rect 119706 248956 119712 249008
rect 119764 248996 119770 249008
rect 119982 248996 119988 249008
rect 119764 248968 119988 248996
rect 119764 248956 119770 248968
rect 119982 248956 119988 248968
rect 120040 248956 120046 249008
rect 156598 248616 156604 248668
rect 156656 248656 156662 248668
rect 212534 248656 212540 248668
rect 156656 248628 212540 248656
rect 156656 248616 156662 248628
rect 212534 248616 212540 248628
rect 212592 248616 212598 248668
rect 68738 248548 68744 248600
rect 68796 248588 68802 248600
rect 126422 248588 126428 248600
rect 68796 248560 126428 248588
rect 68796 248548 68802 248560
rect 126422 248548 126428 248560
rect 126480 248548 126486 248600
rect 159358 248548 159364 248600
rect 159416 248588 159422 248600
rect 218146 248588 218152 248600
rect 159416 248560 218152 248588
rect 159416 248548 159422 248560
rect 218146 248548 218152 248560
rect 218204 248548 218210 248600
rect 119154 248480 119160 248532
rect 119212 248520 119218 248532
rect 119212 248492 162164 248520
rect 119212 248480 119218 248492
rect 162136 248464 162164 248492
rect 69842 248412 69848 248464
rect 69900 248452 69906 248464
rect 126514 248452 126520 248464
rect 69900 248424 126520 248452
rect 69900 248412 69906 248424
rect 126514 248412 126520 248424
rect 126572 248412 126578 248464
rect 162118 248412 162124 248464
rect 162176 248452 162182 248464
rect 223574 248452 223580 248464
rect 162176 248424 223580 248452
rect 162176 248412 162182 248424
rect 223574 248412 223580 248424
rect 223632 248412 223638 248464
rect 121454 248344 121460 248396
rect 121512 248384 121518 248396
rect 121822 248384 121828 248396
rect 121512 248356 121828 248384
rect 121512 248344 121518 248356
rect 121822 248344 121828 248356
rect 121880 248344 121886 248396
rect 119246 247732 119252 247784
rect 119304 247772 119310 247784
rect 127618 247772 127624 247784
rect 119304 247744 127624 247772
rect 119304 247732 119310 247744
rect 127618 247732 127624 247744
rect 127676 247732 127682 247784
rect 10318 247664 10324 247716
rect 10376 247704 10382 247716
rect 67634 247704 67640 247716
rect 10376 247676 67640 247704
rect 10376 247664 10382 247676
rect 67634 247664 67640 247676
rect 67692 247664 67698 247716
rect 119890 247664 119896 247716
rect 119948 247704 119954 247716
rect 172606 247704 172612 247716
rect 119948 247676 172612 247704
rect 119948 247664 119954 247676
rect 172606 247664 172612 247676
rect 172664 247664 172670 247716
rect 127618 247188 127624 247240
rect 127676 247228 127682 247240
rect 200114 247228 200120 247240
rect 127676 247200 200120 247228
rect 127676 247188 127682 247200
rect 200114 247188 200120 247200
rect 200172 247188 200178 247240
rect 133782 247120 133788 247172
rect 133840 247160 133846 247172
rect 213362 247160 213368 247172
rect 133840 247132 213368 247160
rect 133840 247120 133846 247132
rect 213362 247120 213368 247132
rect 213420 247120 213426 247172
rect 121454 247052 121460 247104
rect 121512 247092 121518 247104
rect 230290 247092 230296 247104
rect 121512 247064 230296 247092
rect 121512 247052 121518 247064
rect 230290 247052 230296 247064
rect 230348 247052 230354 247104
rect 121362 246440 121368 246492
rect 121420 246480 121426 246492
rect 173894 246480 173900 246492
rect 121420 246452 173900 246480
rect 121420 246440 121426 246452
rect 173894 246440 173900 246452
rect 173952 246440 173958 246492
rect 122190 246372 122196 246424
rect 122248 246412 122254 246424
rect 175458 246412 175464 246424
rect 122248 246384 175464 246412
rect 122248 246372 122254 246384
rect 175458 246372 175464 246384
rect 175516 246372 175522 246424
rect 122006 246304 122012 246356
rect 122064 246344 122070 246356
rect 122374 246344 122380 246356
rect 122064 246316 122380 246344
rect 122064 246304 122070 246316
rect 122374 246304 122380 246316
rect 122432 246344 122438 246356
rect 229462 246344 229468 246356
rect 122432 246316 229468 246344
rect 122432 246304 122438 246316
rect 229462 246304 229468 246316
rect 229520 246304 229526 246356
rect 122650 245692 122656 245744
rect 122708 245732 122714 245744
rect 128998 245732 129004 245744
rect 122708 245704 129004 245732
rect 122708 245692 122714 245704
rect 128998 245692 129004 245704
rect 129056 245692 129062 245744
rect 121454 245624 121460 245676
rect 121512 245664 121518 245676
rect 122006 245664 122012 245676
rect 121512 245636 122012 245664
rect 121512 245624 121518 245636
rect 122006 245624 122012 245636
rect 122064 245664 122070 245676
rect 230198 245664 230204 245676
rect 122064 245636 230204 245664
rect 122064 245624 122070 245636
rect 230198 245624 230204 245636
rect 230256 245624 230262 245676
rect 121270 244944 121276 244996
rect 121328 244984 121334 244996
rect 137278 244984 137284 244996
rect 121328 244956 137284 244984
rect 121328 244944 121334 244956
rect 137278 244944 137284 244956
rect 137336 244944 137342 244996
rect 15838 244876 15844 244928
rect 15896 244916 15902 244928
rect 64506 244916 64512 244928
rect 15896 244888 64512 244916
rect 15896 244876 15902 244888
rect 64506 244876 64512 244888
rect 64564 244876 64570 244928
rect 122098 244876 122104 244928
rect 122156 244916 122162 244928
rect 171134 244916 171140 244928
rect 122156 244888 171140 244916
rect 122156 244876 122162 244888
rect 171134 244876 171140 244888
rect 171192 244876 171198 244928
rect 137278 244468 137284 244520
rect 137336 244508 137342 244520
rect 218054 244508 218060 244520
rect 137336 244480 218060 244508
rect 137336 244468 137342 244480
rect 218054 244468 218060 244480
rect 218112 244468 218118 244520
rect 121454 244400 121460 244452
rect 121512 244440 121518 244452
rect 230934 244440 230940 244452
rect 121512 244412 230940 244440
rect 121512 244400 121518 244412
rect 230934 244400 230940 244412
rect 230992 244400 230998 244452
rect 121638 244332 121644 244384
rect 121696 244372 121702 244384
rect 231302 244372 231308 244384
rect 121696 244344 231308 244372
rect 121696 244332 121702 244344
rect 231302 244332 231308 244344
rect 231360 244332 231366 244384
rect 64506 244264 64512 244316
rect 64564 244304 64570 244316
rect 67634 244304 67640 244316
rect 64564 244276 67640 244304
rect 64564 244264 64570 244276
rect 67634 244264 67640 244276
rect 67692 244264 67698 244316
rect 205634 244264 205640 244316
rect 205692 244304 205698 244316
rect 580166 244304 580172 244316
rect 205692 244276 580172 244304
rect 205692 244264 205698 244276
rect 580166 244264 580172 244276
rect 580224 244264 580230 244316
rect 68186 243584 68192 243636
rect 68244 243624 68250 243636
rect 68830 243624 68836 243636
rect 68244 243596 68836 243624
rect 68244 243584 68250 243596
rect 68830 243584 68836 243596
rect 68888 243584 68894 243636
rect 68370 243516 68376 243568
rect 68428 243556 68434 243568
rect 68646 243556 68652 243568
rect 68428 243528 68652 243556
rect 68428 243516 68434 243528
rect 68646 243516 68652 243528
rect 68704 243516 68710 243568
rect 66990 243448 66996 243500
rect 67048 243488 67054 243500
rect 69474 243488 69480 243500
rect 67048 243460 69480 243488
rect 67048 243448 67054 243460
rect 69474 243448 69480 243460
rect 69532 243448 69538 243500
rect 122282 242972 122288 243024
rect 122340 243012 122346 243024
rect 230106 243012 230112 243024
rect 122340 242984 230112 243012
rect 122340 242972 122346 242984
rect 230106 242972 230112 242984
rect 230164 242972 230170 243024
rect 121546 242904 121552 242956
rect 121604 242944 121610 242956
rect 122098 242944 122104 242956
rect 121604 242916 122104 242944
rect 121604 242904 121610 242916
rect 122098 242904 122104 242916
rect 122156 242944 122162 242956
rect 231946 242944 231952 242956
rect 122156 242916 231952 242944
rect 122156 242904 122162 242916
rect 231946 242904 231952 242916
rect 232004 242904 232010 242956
rect 168282 242156 168288 242208
rect 168340 242196 168346 242208
rect 205634 242196 205640 242208
rect 168340 242168 205640 242196
rect 168340 242156 168346 242168
rect 205634 242156 205640 242168
rect 205692 242156 205698 242208
rect 121546 241544 121552 241596
rect 121604 241584 121610 241596
rect 230014 241584 230020 241596
rect 121604 241556 230020 241584
rect 121604 241544 121610 241556
rect 230014 241544 230020 241556
rect 230072 241544 230078 241596
rect 121454 241476 121460 241528
rect 121512 241516 121518 241528
rect 231026 241516 231032 241528
rect 121512 241488 231032 241516
rect 121512 241476 121518 241488
rect 231026 241476 231032 241488
rect 231084 241476 231090 241528
rect 67082 240932 67088 240984
rect 67140 240972 67146 240984
rect 68370 240972 68376 240984
rect 67140 240944 68376 240972
rect 67140 240932 67146 240944
rect 68370 240932 68376 240944
rect 68428 240932 68434 240984
rect 125134 240728 125140 240780
rect 125192 240768 125198 240780
rect 159450 240768 159456 240780
rect 125192 240740 159456 240768
rect 125192 240728 125198 240740
rect 159450 240728 159456 240740
rect 159508 240728 159514 240780
rect 177298 240728 177304 240780
rect 177356 240768 177362 240780
rect 208946 240768 208952 240780
rect 177356 240740 208952 240768
rect 177356 240728 177362 240740
rect 208946 240728 208952 240740
rect 209004 240728 209010 240780
rect 3050 240116 3056 240168
rect 3108 240156 3114 240168
rect 66898 240156 66904 240168
rect 3108 240128 66904 240156
rect 3108 240116 3114 240128
rect 66898 240116 66904 240128
rect 66956 240116 66962 240168
rect 159450 240116 159456 240168
rect 159508 240156 159514 240168
rect 207658 240156 207664 240168
rect 159508 240128 207664 240156
rect 159508 240116 159514 240128
rect 207658 240116 207664 240128
rect 207716 240116 207722 240168
rect 121822 239436 121828 239488
rect 121880 239476 121886 239488
rect 147582 239476 147588 239488
rect 121880 239448 147588 239476
rect 121880 239436 121886 239448
rect 147582 239436 147588 239448
rect 147640 239436 147646 239488
rect 124122 239368 124128 239420
rect 124180 239408 124186 239420
rect 158070 239408 158076 239420
rect 124180 239380 158076 239408
rect 124180 239368 124186 239380
rect 158070 239368 158076 239380
rect 158128 239368 158134 239420
rect 168926 239368 168932 239420
rect 168984 239408 168990 239420
rect 282914 239408 282920 239420
rect 168984 239380 282920 239408
rect 168984 239368 168990 239380
rect 282914 239368 282920 239380
rect 282972 239368 282978 239420
rect 158070 238824 158076 238876
rect 158128 238864 158134 238876
rect 190638 238864 190644 238876
rect 158128 238836 190644 238864
rect 158128 238824 158134 238836
rect 190638 238824 190644 238836
rect 190696 238824 190702 238876
rect 147582 238756 147588 238808
rect 147640 238796 147646 238808
rect 231210 238796 231216 238808
rect 147640 238768 231216 238796
rect 147640 238756 147646 238768
rect 231210 238756 231216 238768
rect 231268 238756 231274 238808
rect 127802 237532 127808 237584
rect 127860 237572 127866 237584
rect 131942 237572 131948 237584
rect 127860 237544 131948 237572
rect 127860 237532 127866 237544
rect 131942 237532 131948 237544
rect 132000 237572 132006 237584
rect 202874 237572 202880 237584
rect 132000 237544 202880 237572
rect 132000 237532 132006 237544
rect 202874 237532 202880 237544
rect 202932 237532 202938 237584
rect 121822 237464 121828 237516
rect 121880 237504 121886 237516
rect 230750 237504 230756 237516
rect 121880 237476 230756 237504
rect 121880 237464 121886 237476
rect 230750 237464 230756 237476
rect 230808 237464 230814 237516
rect 231118 237436 231124 237448
rect 122806 237408 231124 237436
rect 121362 237328 121368 237380
rect 121420 237368 121426 237380
rect 122806 237368 122834 237408
rect 231118 237396 231124 237408
rect 231176 237396 231182 237448
rect 121420 237340 122834 237368
rect 121420 237328 121426 237340
rect 130378 236784 130384 236836
rect 130436 236824 130442 236836
rect 177114 236824 177120 236836
rect 130436 236796 177120 236824
rect 130436 236784 130442 236796
rect 177114 236784 177120 236796
rect 177172 236784 177178 236836
rect 186130 236784 186136 236836
rect 186188 236824 186194 236836
rect 195238 236824 195244 236836
rect 186188 236796 195244 236824
rect 186188 236784 186194 236796
rect 195238 236784 195244 236796
rect 195296 236784 195302 236836
rect 128998 236716 129004 236768
rect 129056 236756 129062 236768
rect 232682 236756 232688 236768
rect 129056 236728 232688 236756
rect 129056 236716 129062 236728
rect 232682 236716 232688 236728
rect 232740 236716 232746 236768
rect 169110 236648 169116 236700
rect 169168 236688 169174 236700
rect 580350 236688 580356 236700
rect 169168 236660 580356 236688
rect 169168 236648 169174 236660
rect 580350 236648 580356 236660
rect 580408 236648 580414 236700
rect 122742 235968 122748 236020
rect 122800 236008 122806 236020
rect 230566 236008 230572 236020
rect 122800 235980 230572 236008
rect 122800 235968 122806 235980
rect 230566 235968 230572 235980
rect 230624 235968 230630 236020
rect 126698 234744 126704 234796
rect 126756 234784 126762 234796
rect 133230 234784 133236 234796
rect 126756 234756 133236 234784
rect 126756 234744 126762 234756
rect 133230 234744 133236 234756
rect 133288 234784 133294 234796
rect 226702 234784 226708 234796
rect 133288 234756 226708 234784
rect 133288 234744 133294 234756
rect 226702 234744 226708 234756
rect 226760 234744 226766 234796
rect 122282 234676 122288 234728
rect 122340 234716 122346 234728
rect 229554 234716 229560 234728
rect 122340 234688 229560 234716
rect 122340 234676 122346 234688
rect 229554 234676 229560 234688
rect 229612 234676 229618 234728
rect 122466 234608 122472 234660
rect 122524 234648 122530 234660
rect 230474 234648 230480 234660
rect 122524 234620 230480 234648
rect 122524 234608 122530 234620
rect 230474 234608 230480 234620
rect 230532 234608 230538 234660
rect 190454 233928 190460 233980
rect 190512 233968 190518 233980
rect 191006 233968 191012 233980
rect 190512 233940 191012 233968
rect 190512 233928 190518 233940
rect 191006 233928 191012 233940
rect 191064 233928 191070 233980
rect 194594 233928 194600 233980
rect 194652 233968 194658 233980
rect 195422 233968 195428 233980
rect 194652 233940 195428 233968
rect 194652 233928 194658 233940
rect 195422 233928 195428 233940
rect 195480 233928 195486 233980
rect 218054 233928 218060 233980
rect 218112 233968 218118 233980
rect 218606 233968 218612 233980
rect 218112 233940 218612 233968
rect 218112 233928 218118 233940
rect 218606 233928 218612 233940
rect 218664 233928 218670 233980
rect 68462 233860 68468 233912
rect 68520 233900 68526 233912
rect 68738 233900 68744 233912
rect 68520 233872 68744 233900
rect 68520 233860 68526 233872
rect 68738 233860 68744 233872
rect 68796 233860 68802 233912
rect 126606 233860 126612 233912
rect 126664 233900 126670 233912
rect 229278 233900 229284 233912
rect 126664 233872 229284 233900
rect 126664 233860 126670 233872
rect 229278 233860 229284 233872
rect 229336 233860 229342 233912
rect 122466 233248 122472 233300
rect 122524 233288 122530 233300
rect 230382 233288 230388 233300
rect 122524 233260 230388 233288
rect 122524 233248 122530 233260
rect 230382 233248 230388 233260
rect 230440 233248 230446 233300
rect 121270 233180 121276 233232
rect 121328 233220 121334 233232
rect 122006 233220 122012 233232
rect 121328 233192 122012 233220
rect 121328 233180 121334 233192
rect 122006 233180 122012 233192
rect 122064 233180 122070 233232
rect 186130 233220 186136 233232
rect 122116 233192 186136 233220
rect 121086 233112 121092 233164
rect 121144 233152 121150 233164
rect 122116 233152 122144 233192
rect 186130 233180 186136 233192
rect 186188 233180 186194 233232
rect 215938 233180 215944 233232
rect 215996 233220 216002 233232
rect 217042 233220 217048 233232
rect 215996 233192 217048 233220
rect 215996 233180 216002 233192
rect 217042 233180 217048 233192
rect 217100 233180 217106 233232
rect 331214 233220 331220 233232
rect 219406 233192 331220 233220
rect 171226 233152 171232 233164
rect 121144 233124 122144 233152
rect 122806 233124 171232 233152
rect 121144 233112 121150 233124
rect 119338 233044 119344 233096
rect 119396 233084 119402 233096
rect 122806 233084 122834 233124
rect 171226 233112 171232 233124
rect 171284 233152 171290 233164
rect 180058 233152 180064 233164
rect 171284 233124 180064 233152
rect 171284 233112 171290 233124
rect 180058 233112 180064 233124
rect 180116 233112 180122 233164
rect 210418 233112 210424 233164
rect 210476 233152 210482 233164
rect 214466 233152 214472 233164
rect 210476 233124 214472 233152
rect 210476 233112 210482 233124
rect 214466 233112 214472 233124
rect 214524 233112 214530 233164
rect 119396 233056 122834 233084
rect 119396 233044 119402 233056
rect 213362 233044 213368 233096
rect 213420 233084 213426 233096
rect 219406 233084 219434 233192
rect 331214 233180 331220 233192
rect 331272 233180 331278 233232
rect 222838 233112 222844 233164
rect 222896 233152 222902 233164
rect 226058 233152 226064 233164
rect 222896 233124 226064 233152
rect 222896 233112 222902 233124
rect 226058 233112 226064 233124
rect 226116 233112 226122 233164
rect 213420 233056 219434 233084
rect 213420 233044 213426 233056
rect 121178 232772 121184 232824
rect 121236 232812 121242 232824
rect 134610 232812 134616 232824
rect 121236 232784 134616 232812
rect 121236 232772 121242 232784
rect 134610 232772 134616 232784
rect 134668 232772 134674 232824
rect 119706 232704 119712 232756
rect 119764 232744 119770 232756
rect 138658 232744 138664 232756
rect 119764 232716 138664 232744
rect 119764 232704 119770 232716
rect 138658 232704 138664 232716
rect 138716 232704 138722 232756
rect 120994 232636 121000 232688
rect 121052 232676 121058 232688
rect 166810 232676 166816 232688
rect 121052 232648 166816 232676
rect 121052 232636 121058 232648
rect 166810 232636 166816 232648
rect 166868 232636 166874 232688
rect 189350 232676 189356 232688
rect 180766 232648 189356 232676
rect 66622 232568 66628 232620
rect 66680 232608 66686 232620
rect 68738 232608 68744 232620
rect 66680 232580 68744 232608
rect 66680 232568 66686 232580
rect 68738 232568 68744 232580
rect 68796 232568 68802 232620
rect 133322 232568 133328 232620
rect 133380 232608 133386 232620
rect 180766 232608 180794 232648
rect 189350 232636 189356 232648
rect 189408 232636 189414 232688
rect 133380 232580 180794 232608
rect 133380 232568 133386 232580
rect 181438 232568 181444 232620
rect 181496 232608 181502 232620
rect 181496 232580 190454 232608
rect 181496 232568 181502 232580
rect 119798 232500 119804 232552
rect 119856 232540 119862 232552
rect 181622 232540 181628 232552
rect 119856 232512 181628 232540
rect 119856 232500 119862 232512
rect 181622 232500 181628 232512
rect 181680 232500 181686 232552
rect 190426 232540 190454 232580
rect 198366 232540 198372 232552
rect 190426 232512 198372 232540
rect 198366 232500 198372 232512
rect 198424 232500 198430 232552
rect 226058 232500 226064 232552
rect 226116 232540 226122 232552
rect 412634 232540 412640 232552
rect 226116 232512 412640 232540
rect 226116 232500 226122 232512
rect 412634 232500 412640 232512
rect 412692 232500 412698 232552
rect 166902 232092 166908 232144
rect 166960 232132 166966 232144
rect 215754 232132 215760 232144
rect 166960 232104 215760 232132
rect 166960 232092 166966 232104
rect 215754 232092 215760 232104
rect 215812 232092 215818 232144
rect 140774 232024 140780 232076
rect 140832 232064 140838 232076
rect 141418 232064 141424 232076
rect 140832 232036 141424 232064
rect 140832 232024 140838 232036
rect 141418 232024 141424 232036
rect 141476 232064 141482 232076
rect 192570 232064 192576 232076
rect 141476 232036 192576 232064
rect 141476 232024 141482 232036
rect 192570 232024 192576 232036
rect 192628 232024 192634 232076
rect 204898 232024 204904 232076
rect 204956 232064 204962 232076
rect 234614 232064 234620 232076
rect 204956 232036 234620 232064
rect 204956 232024 204962 232036
rect 234614 232024 234620 232036
rect 234672 232024 234678 232076
rect 166810 231956 166816 232008
rect 166868 231996 166874 232008
rect 221550 231996 221556 232008
rect 166868 231968 221556 231996
rect 166868 231956 166874 231968
rect 221550 231956 221556 231968
rect 221608 231956 221614 232008
rect 223482 231956 223488 232008
rect 223540 231996 223546 232008
rect 233234 231996 233240 232008
rect 223540 231968 233240 231996
rect 223540 231956 223546 231968
rect 233234 231956 233240 231968
rect 233292 231956 233298 232008
rect 134610 231888 134616 231940
rect 134668 231928 134674 231940
rect 206094 231928 206100 231940
rect 134668 231900 206100 231928
rect 134668 231888 134674 231900
rect 206094 231888 206100 231900
rect 206152 231888 206158 231940
rect 138658 231820 138664 231872
rect 138716 231860 138722 231872
rect 210602 231860 210608 231872
rect 138716 231832 210608 231860
rect 138716 231820 138722 231832
rect 210602 231820 210608 231832
rect 210660 231820 210666 231872
rect 222194 231820 222200 231872
rect 222252 231860 222258 231872
rect 234706 231860 234712 231872
rect 222252 231832 234712 231860
rect 222252 231820 222258 231832
rect 234706 231820 234712 231832
rect 234764 231820 234770 231872
rect 173986 231208 173992 231260
rect 174044 231248 174050 231260
rect 175182 231248 175188 231260
rect 174044 231220 175188 231248
rect 174044 231208 174050 231220
rect 175182 231208 175188 231220
rect 175240 231208 175246 231260
rect 126514 231072 126520 231124
rect 126572 231112 126578 231124
rect 150434 231112 150440 231124
rect 126572 231084 150440 231112
rect 126572 231072 126578 231084
rect 150434 231072 150440 231084
rect 150492 231072 150498 231124
rect 168190 231072 168196 231124
rect 168248 231112 168254 231124
rect 579982 231112 579988 231124
rect 168248 231084 579988 231112
rect 168248 231072 168254 231084
rect 579982 231072 579988 231084
rect 580040 231072 580046 231124
rect 121730 230868 121736 230920
rect 121788 230908 121794 230920
rect 122282 230908 122288 230920
rect 121788 230880 122288 230908
rect 121788 230868 121794 230880
rect 122282 230868 122288 230880
rect 122340 230908 122346 230920
rect 229094 230908 229100 230920
rect 122340 230880 229100 230908
rect 122340 230868 122346 230880
rect 229094 230868 229100 230880
rect 229152 230868 229158 230920
rect 121454 230800 121460 230852
rect 121512 230840 121518 230852
rect 230658 230840 230664 230852
rect 121512 230812 230664 230840
rect 121512 230800 121518 230812
rect 230658 230800 230664 230812
rect 230716 230800 230722 230852
rect 169294 230732 169300 230784
rect 169352 230772 169358 230784
rect 179414 230772 179420 230784
rect 169352 230744 179420 230772
rect 169352 230732 169358 230744
rect 179414 230732 179420 230744
rect 179472 230732 179478 230784
rect 169202 230664 169208 230716
rect 169260 230704 169266 230716
rect 182450 230704 182456 230716
rect 169260 230676 182456 230704
rect 169260 230664 169266 230676
rect 182450 230664 182456 230676
rect 182508 230664 182514 230716
rect 150434 230596 150440 230648
rect 150492 230636 150498 230648
rect 150492 230608 161474 230636
rect 150492 230596 150498 230608
rect 65794 230460 65800 230512
rect 65852 230500 65858 230512
rect 67634 230500 67640 230512
rect 65852 230472 67640 230500
rect 65852 230460 65858 230472
rect 67634 230460 67640 230472
rect 67692 230460 67698 230512
rect 161446 230500 161474 230608
rect 170030 230596 170036 230648
rect 170088 230636 170094 230648
rect 183554 230636 183560 230648
rect 170088 230608 183560 230636
rect 170088 230596 170094 230608
rect 183554 230596 183560 230608
rect 183612 230636 183618 230648
rect 184842 230636 184848 230648
rect 183612 230608 184848 230636
rect 183612 230596 183618 230608
rect 184842 230596 184848 230608
rect 184900 230596 184906 230648
rect 198366 230596 198372 230648
rect 198424 230636 198430 230648
rect 235350 230636 235356 230648
rect 198424 230608 235356 230636
rect 198424 230596 198430 230608
rect 235350 230596 235356 230608
rect 235408 230596 235414 230648
rect 169386 230528 169392 230580
rect 169444 230568 169450 230580
rect 173986 230568 173992 230580
rect 169444 230540 173992 230568
rect 169444 230528 169450 230540
rect 173986 230528 173992 230540
rect 174044 230528 174050 230580
rect 161446 230472 167776 230500
rect 65886 230392 65892 230444
rect 65944 230432 65950 230444
rect 67726 230432 67732 230444
rect 65944 230404 67732 230432
rect 65944 230392 65950 230404
rect 67726 230392 67732 230404
rect 67784 230392 67790 230444
rect 167748 230432 167776 230472
rect 169478 230460 169484 230512
rect 169536 230500 169542 230512
rect 171134 230500 171140 230512
rect 169536 230472 171140 230500
rect 169536 230460 169542 230472
rect 171134 230460 171140 230472
rect 171192 230460 171198 230512
rect 170674 230432 170680 230444
rect 167748 230404 170680 230432
rect 170674 230392 170680 230404
rect 170732 230432 170738 230444
rect 173158 230432 173164 230444
rect 170732 230404 173164 230432
rect 170732 230392 170738 230404
rect 173158 230392 173164 230404
rect 173216 230392 173222 230444
rect 229922 230392 229928 230444
rect 229980 230432 229986 230444
rect 231946 230432 231952 230444
rect 229980 230404 231952 230432
rect 229980 230392 229986 230404
rect 231946 230392 231952 230404
rect 232004 230392 232010 230444
rect 163498 229848 163504 229900
rect 163556 229888 163562 229900
rect 232314 229888 232320 229900
rect 163556 229860 232320 229888
rect 163556 229848 163562 229860
rect 232314 229848 232320 229860
rect 232372 229848 232378 229900
rect 120902 229780 120908 229832
rect 120960 229820 120966 229832
rect 166994 229820 167000 229832
rect 120960 229792 167000 229820
rect 120960 229780 120966 229792
rect 166994 229780 167000 229792
rect 167052 229780 167058 229832
rect 166258 229712 166264 229764
rect 166316 229752 166322 229764
rect 231946 229752 231952 229764
rect 166316 229724 231952 229752
rect 166316 229712 166322 229724
rect 231946 229712 231952 229724
rect 232004 229712 232010 229764
rect 166350 229644 166356 229696
rect 166408 229684 166414 229696
rect 232130 229684 232136 229696
rect 166408 229656 232136 229684
rect 166408 229644 166414 229656
rect 232130 229644 232136 229656
rect 232188 229644 232194 229696
rect 166442 229576 166448 229628
rect 166500 229616 166506 229628
rect 232222 229616 232228 229628
rect 166500 229588 232228 229616
rect 166500 229576 166506 229588
rect 232222 229576 232228 229588
rect 232280 229576 232286 229628
rect 166718 229508 166724 229560
rect 166776 229548 166782 229560
rect 232498 229548 232504 229560
rect 166776 229520 232504 229548
rect 166776 229508 166782 229520
rect 232498 229508 232504 229520
rect 232556 229508 232562 229560
rect 166534 229440 166540 229492
rect 166592 229480 166598 229492
rect 232406 229480 232412 229492
rect 166592 229452 232412 229480
rect 166592 229440 166598 229452
rect 232406 229440 232412 229452
rect 232464 229440 232470 229492
rect 165430 229372 165436 229424
rect 165488 229412 165494 229424
rect 232590 229412 232596 229424
rect 165488 229384 232596 229412
rect 165488 229372 165494 229384
rect 232590 229372 232596 229384
rect 232648 229372 232654 229424
rect 162394 229304 162400 229356
rect 162452 229344 162458 229356
rect 232038 229344 232044 229356
rect 162452 229316 232044 229344
rect 162452 229304 162458 229316
rect 232038 229304 232044 229316
rect 232096 229304 232102 229356
rect 144270 229168 144276 229220
rect 144328 229208 144334 229220
rect 231854 229208 231860 229220
rect 144328 229180 231860 229208
rect 144328 229168 144334 229180
rect 231854 229168 231860 229180
rect 231912 229168 231918 229220
rect 121454 229100 121460 229152
rect 121512 229140 121518 229152
rect 229278 229140 229284 229152
rect 121512 229112 229284 229140
rect 121512 229100 121518 229112
rect 229278 229100 229284 229112
rect 229336 229100 229342 229152
rect 229370 229100 229376 229152
rect 229428 229140 229434 229152
rect 230842 229140 230848 229152
rect 229428 229112 230848 229140
rect 229428 229100 229434 229112
rect 230842 229100 230848 229112
rect 230900 229100 230906 229152
rect 125042 229032 125048 229084
rect 125100 229072 125106 229084
rect 167086 229072 167092 229084
rect 125100 229044 167092 229072
rect 125100 229032 125106 229044
rect 167086 229032 167092 229044
rect 167144 229032 167150 229084
rect 231026 229032 231032 229084
rect 231084 229072 231090 229084
rect 231394 229072 231400 229084
rect 231084 229044 231400 229072
rect 231084 229032 231090 229044
rect 231394 229032 231400 229044
rect 231452 229072 231458 229084
rect 233970 229072 233976 229084
rect 231452 229044 233976 229072
rect 231452 229032 231458 229044
rect 233970 229032 233976 229044
rect 234028 229032 234034 229084
rect 164878 226312 164884 226364
rect 164936 226352 164942 226364
rect 167546 226352 167552 226364
rect 164936 226324 167552 226352
rect 164936 226312 164942 226324
rect 167546 226312 167552 226324
rect 167604 226312 167610 226364
rect 229646 226312 229652 226364
rect 229704 226352 229710 226364
rect 548610 226352 548616 226364
rect 229704 226324 548616 226352
rect 229704 226312 229710 226324
rect 548610 226312 548616 226324
rect 548668 226312 548674 226364
rect 63494 225564 63500 225616
rect 63552 225604 63558 225616
rect 64598 225604 64604 225616
rect 63552 225576 64604 225604
rect 63552 225564 63558 225576
rect 64598 225564 64604 225576
rect 64656 225604 64662 225616
rect 67818 225604 67824 225616
rect 64656 225576 67824 225604
rect 64656 225564 64662 225576
rect 67818 225564 67824 225576
rect 67876 225564 67882 225616
rect 122466 225564 122472 225616
rect 122524 225604 122530 225616
rect 165430 225604 165436 225616
rect 122524 225576 165436 225604
rect 122524 225564 122530 225576
rect 165430 225564 165436 225576
rect 165488 225564 165494 225616
rect 66898 225292 66904 225344
rect 66956 225332 66962 225344
rect 68738 225332 68744 225344
rect 66956 225304 68744 225332
rect 66956 225292 66962 225304
rect 68738 225292 68744 225304
rect 68796 225292 68802 225344
rect 15838 224952 15844 225004
rect 15896 224992 15902 225004
rect 63494 224992 63500 225004
rect 15896 224964 63500 224992
rect 15896 224952 15902 224964
rect 63494 224952 63500 224964
rect 63552 224952 63558 225004
rect 119890 224952 119896 225004
rect 119948 224992 119954 225004
rect 121546 224992 121552 225004
rect 119948 224964 121552 224992
rect 119948 224952 119954 224964
rect 121546 224952 121552 224964
rect 121604 224952 121610 225004
rect 139394 224952 139400 225004
rect 139452 224992 139458 225004
rect 167086 224992 167092 225004
rect 139452 224964 167092 224992
rect 139452 224952 139458 224964
rect 167086 224952 167092 224964
rect 167144 224952 167150 225004
rect 121454 224884 121460 224936
rect 121512 224924 121518 224936
rect 166718 224924 166724 224936
rect 121512 224896 166724 224924
rect 121512 224884 121518 224896
rect 166718 224884 166724 224896
rect 166776 224884 166782 224936
rect 124030 224816 124036 224868
rect 124088 224856 124094 224868
rect 167086 224856 167092 224868
rect 124088 224828 167092 224856
rect 124088 224816 124094 224828
rect 167086 224816 167092 224828
rect 167144 224816 167150 224868
rect 230934 223524 230940 223576
rect 230992 223564 230998 223576
rect 558914 223564 558920 223576
rect 230992 223536 558920 223564
rect 230992 223524 230998 223536
rect 558914 223524 558920 223536
rect 558972 223524 558978 223576
rect 125042 222164 125048 222216
rect 125100 222204 125106 222216
rect 167086 222204 167092 222216
rect 125100 222176 167092 222204
rect 125100 222164 125106 222176
rect 167086 222164 167092 222176
rect 167144 222164 167150 222216
rect 121454 222028 121460 222080
rect 121512 222068 121518 222080
rect 123662 222068 123668 222080
rect 121512 222040 123668 222068
rect 121512 222028 121518 222040
rect 123662 222028 123668 222040
rect 123720 222028 123726 222080
rect 124950 221416 124956 221468
rect 125008 221456 125014 221468
rect 167454 221456 167460 221468
rect 125008 221428 167460 221456
rect 125008 221416 125014 221428
rect 167454 221416 167460 221428
rect 167512 221416 167518 221468
rect 65610 220804 65616 220856
rect 65668 220844 65674 220856
rect 68002 220844 68008 220856
rect 65668 220816 68008 220844
rect 65668 220804 65674 220816
rect 68002 220804 68008 220816
rect 68060 220804 68066 220856
rect 120442 220736 120448 220788
rect 120500 220776 120506 220788
rect 166534 220776 166540 220788
rect 120500 220748 166540 220776
rect 120500 220736 120506 220748
rect 166534 220736 166540 220748
rect 166592 220736 166598 220788
rect 67450 219444 67456 219496
rect 67508 219484 67514 219496
rect 68922 219484 68928 219496
rect 67508 219456 68928 219484
rect 67508 219444 67514 219456
rect 68922 219444 68928 219456
rect 68980 219444 68986 219496
rect 119522 219376 119528 219428
rect 119580 219416 119586 219428
rect 163498 219416 163504 219428
rect 119580 219388 163504 219416
rect 119580 219376 119586 219388
rect 163498 219376 163504 219388
rect 163556 219376 163562 219428
rect 235350 219376 235356 219428
rect 235408 219416 235414 219428
rect 580166 219416 580172 219428
rect 235408 219388 580172 219416
rect 235408 219376 235414 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 153838 219308 153844 219360
rect 153896 219348 153902 219360
rect 167086 219348 167092 219360
rect 153896 219320 167092 219348
rect 153896 219308 153902 219320
rect 167086 219308 167092 219320
rect 167144 219308 167150 219360
rect 119154 218424 119160 218476
rect 119212 218464 119218 218476
rect 119522 218464 119528 218476
rect 119212 218436 119528 218464
rect 119212 218424 119218 218436
rect 119522 218424 119528 218436
rect 119580 218424 119586 218476
rect 120718 218084 120724 218136
rect 120776 218124 120782 218136
rect 121546 218124 121552 218136
rect 120776 218096 121552 218124
rect 120776 218084 120782 218096
rect 121546 218084 121552 218096
rect 121604 218084 121610 218136
rect 65886 218016 65892 218068
rect 65944 218056 65950 218068
rect 68186 218056 68192 218068
rect 65944 218028 68192 218056
rect 65944 218016 65950 218028
rect 68186 218016 68192 218028
rect 68244 218016 68250 218068
rect 120994 218016 121000 218068
rect 121052 218056 121058 218068
rect 121454 218056 121460 218068
rect 121052 218028 121460 218056
rect 121052 218016 121058 218028
rect 121454 218016 121460 218028
rect 121512 218016 121518 218068
rect 119430 217948 119436 218000
rect 119488 217988 119494 218000
rect 167086 217988 167092 218000
rect 119488 217960 167092 217988
rect 119488 217948 119494 217960
rect 167086 217948 167092 217960
rect 167144 217948 167150 218000
rect 232682 217948 232688 218000
rect 232740 217988 232746 218000
rect 233878 217988 233884 218000
rect 232740 217960 233884 217988
rect 232740 217948 232746 217960
rect 233878 217948 233884 217960
rect 233936 217948 233942 218000
rect 122006 217268 122012 217320
rect 122064 217308 122070 217320
rect 166442 217308 166448 217320
rect 122064 217280 166448 217308
rect 122064 217268 122070 217280
rect 166442 217268 166448 217280
rect 166500 217268 166506 217320
rect 66806 216656 66812 216708
rect 66864 216696 66870 216708
rect 68370 216696 68376 216708
rect 66864 216668 68376 216696
rect 66864 216656 66870 216668
rect 68370 216656 68376 216668
rect 68428 216656 68434 216708
rect 121454 215976 121460 216028
rect 121512 216016 121518 216028
rect 148410 216016 148416 216028
rect 121512 215988 148416 216016
rect 121512 215976 121518 215988
rect 148410 215976 148416 215988
rect 148468 215976 148474 216028
rect 123754 215908 123760 215960
rect 123812 215948 123818 215960
rect 162854 215948 162860 215960
rect 123812 215920 162860 215948
rect 123812 215908 123818 215920
rect 162854 215908 162860 215920
rect 162912 215948 162918 215960
rect 167086 215948 167092 215960
rect 162912 215920 167092 215948
rect 162912 215908 162918 215920
rect 167086 215908 167092 215920
rect 167144 215908 167150 215960
rect 64414 215296 64420 215348
rect 64472 215336 64478 215348
rect 67634 215336 67640 215348
rect 64472 215308 67640 215336
rect 64472 215296 64478 215308
rect 67634 215296 67640 215308
rect 67692 215296 67698 215348
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 15838 215268 15844 215280
rect 3384 215240 15844 215268
rect 3384 215228 3390 215240
rect 15838 215228 15844 215240
rect 15896 215228 15902 215280
rect 123938 214616 123944 214668
rect 123996 214656 124002 214668
rect 144914 214656 144920 214668
rect 123996 214628 144920 214656
rect 123996 214616 124002 214628
rect 144914 214616 144920 214628
rect 144972 214656 144978 214668
rect 145926 214656 145932 214668
rect 144972 214628 145932 214656
rect 144972 214616 144978 214628
rect 145926 214616 145932 214628
rect 145984 214616 145990 214668
rect 3786 214548 3792 214600
rect 3844 214588 3850 214600
rect 67634 214588 67640 214600
rect 3844 214560 67640 214588
rect 3844 214548 3850 214560
rect 67634 214548 67640 214560
rect 67692 214548 67698 214600
rect 123846 214548 123852 214600
rect 123904 214588 123910 214600
rect 154574 214588 154580 214600
rect 123904 214560 154580 214588
rect 123904 214548 123910 214560
rect 154574 214548 154580 214560
rect 154632 214588 154638 214600
rect 155678 214588 155684 214600
rect 154632 214560 155684 214588
rect 154632 214548 154638 214560
rect 155678 214548 155684 214560
rect 155736 214548 155742 214600
rect 120810 214004 120816 214056
rect 120868 214044 120874 214056
rect 121546 214044 121552 214056
rect 120868 214016 121552 214044
rect 120868 214004 120874 214016
rect 121546 214004 121552 214016
rect 121604 214004 121610 214056
rect 155678 214004 155684 214056
rect 155736 214044 155742 214056
rect 167178 214044 167184 214056
rect 155736 214016 167184 214044
rect 155736 214004 155742 214016
rect 167178 214004 167184 214016
rect 167236 214004 167242 214056
rect 121454 213936 121460 213988
rect 121512 213976 121518 213988
rect 142982 213976 142988 213988
rect 121512 213948 142988 213976
rect 121512 213936 121518 213948
rect 142982 213936 142988 213948
rect 143040 213936 143046 213988
rect 145926 213936 145932 213988
rect 145984 213976 145990 213988
rect 167086 213976 167092 213988
rect 145984 213948 167092 213976
rect 145984 213936 145990 213948
rect 167086 213936 167092 213948
rect 167144 213936 167150 213988
rect 121730 213868 121736 213920
rect 121788 213908 121794 213920
rect 144270 213908 144276 213920
rect 121788 213880 144276 213908
rect 121788 213868 121794 213880
rect 144270 213868 144276 213880
rect 144328 213868 144334 213920
rect 119982 212848 119988 212900
rect 120040 212888 120046 212900
rect 122098 212888 122104 212900
rect 120040 212860 122104 212888
rect 120040 212848 120046 212860
rect 122098 212848 122104 212860
rect 122156 212848 122162 212900
rect 121914 212508 121920 212560
rect 121972 212548 121978 212560
rect 156782 212548 156788 212560
rect 121972 212520 156788 212548
rect 121972 212508 121978 212520
rect 156782 212508 156788 212520
rect 156840 212508 156846 212560
rect 121178 212440 121184 212492
rect 121236 212480 121242 212492
rect 122466 212480 122472 212492
rect 121236 212452 122472 212480
rect 121236 212440 121242 212452
rect 122466 212440 122472 212452
rect 122524 212440 122530 212492
rect 121454 211760 121460 211812
rect 121512 211800 121518 211812
rect 122006 211800 122012 211812
rect 121512 211772 122012 211800
rect 121512 211760 121518 211772
rect 122006 211760 122012 211772
rect 122064 211800 122070 211812
rect 166350 211800 166356 211812
rect 122064 211772 166356 211800
rect 122064 211760 122070 211772
rect 166350 211760 166356 211772
rect 166408 211760 166414 211812
rect 121454 211624 121460 211676
rect 121512 211664 121518 211676
rect 121914 211664 121920 211676
rect 121512 211636 121920 211664
rect 121512 211624 121518 211636
rect 121914 211624 121920 211636
rect 121972 211624 121978 211676
rect 162210 211488 162216 211540
rect 162268 211528 162274 211540
rect 167086 211528 167092 211540
rect 162268 211500 167092 211528
rect 162268 211488 162274 211500
rect 167086 211488 167092 211500
rect 167144 211488 167150 211540
rect 162302 210808 162308 210860
rect 162360 210848 162366 210860
rect 167086 210848 167092 210860
rect 162360 210820 167092 210848
rect 162360 210808 162366 210820
rect 167086 210808 167092 210820
rect 167144 210808 167150 210860
rect 123570 209720 123576 209772
rect 123628 209760 123634 209772
rect 168190 209760 168196 209772
rect 123628 209732 168196 209760
rect 123628 209720 123634 209732
rect 168190 209720 168196 209732
rect 168248 209720 168254 209772
rect 230382 209720 230388 209772
rect 230440 209760 230446 209772
rect 234062 209760 234068 209772
rect 230440 209732 234068 209760
rect 230440 209720 230446 209732
rect 234062 209720 234068 209732
rect 234120 209720 234126 209772
rect 229830 208360 229836 208412
rect 229888 208400 229894 208412
rect 230382 208400 230388 208412
rect 229888 208372 230388 208400
rect 229888 208360 229894 208372
rect 230382 208360 230388 208372
rect 230440 208360 230446 208412
rect 124858 207612 124864 207664
rect 124916 207652 124922 207664
rect 158714 207652 158720 207664
rect 124916 207624 158720 207652
rect 124916 207612 124922 207624
rect 158714 207612 158720 207624
rect 158772 207612 158778 207664
rect 158714 207000 158720 207052
rect 158772 207040 158778 207052
rect 167086 207040 167092 207052
rect 158772 207012 167092 207040
rect 158772 207000 158778 207012
rect 167086 207000 167092 207012
rect 167144 207000 167150 207052
rect 548610 206932 548616 206984
rect 548668 206972 548674 206984
rect 579982 206972 579988 206984
rect 548668 206944 579988 206972
rect 548668 206932 548674 206944
rect 579982 206932 579988 206944
rect 580040 206932 580046 206984
rect 137922 206388 137928 206440
rect 137980 206428 137986 206440
rect 167086 206428 167092 206440
rect 137980 206400 167092 206428
rect 137980 206388 137986 206400
rect 167086 206388 167092 206400
rect 167144 206388 167150 206440
rect 121546 206320 121552 206372
rect 121604 206360 121610 206372
rect 122098 206360 122104 206372
rect 121604 206332 122104 206360
rect 121604 206320 121610 206332
rect 122098 206320 122104 206332
rect 122156 206360 122162 206372
rect 162394 206360 162400 206372
rect 122156 206332 162400 206360
rect 122156 206320 122162 206332
rect 162394 206320 162400 206332
rect 162452 206320 162458 206372
rect 123478 206252 123484 206304
rect 123536 206292 123542 206304
rect 167086 206292 167092 206304
rect 123536 206264 167092 206292
rect 123536 206252 123542 206264
rect 167086 206252 167092 206264
rect 167144 206252 167150 206304
rect 67358 205640 67364 205692
rect 67416 205680 67422 205692
rect 68370 205680 68376 205692
rect 67416 205652 68376 205680
rect 67416 205640 67422 205652
rect 68370 205640 68376 205652
rect 68428 205640 68434 205692
rect 121086 205640 121092 205692
rect 121144 205680 121150 205692
rect 122282 205680 122288 205692
rect 121144 205652 122288 205680
rect 121144 205640 121150 205652
rect 122282 205640 122288 205652
rect 122340 205640 122346 205692
rect 232682 205640 232688 205692
rect 232740 205680 232746 205692
rect 548518 205680 548524 205692
rect 232740 205652 548524 205680
rect 232740 205640 232746 205652
rect 548518 205640 548524 205652
rect 548576 205640 548582 205692
rect 11698 205572 11704 205624
rect 11756 205612 11762 205624
rect 67818 205612 67824 205624
rect 11756 205584 67824 205612
rect 11756 205572 11762 205584
rect 67818 205572 67824 205584
rect 67876 205572 67882 205624
rect 68002 204892 68008 204944
rect 68060 204932 68066 204944
rect 69382 204932 69388 204944
rect 68060 204904 69388 204932
rect 68060 204892 68066 204904
rect 69382 204892 69388 204904
rect 69440 204892 69446 204944
rect 122558 204892 122564 204944
rect 122616 204932 122622 204944
rect 166258 204932 166264 204944
rect 122616 204904 166264 204932
rect 122616 204892 122622 204904
rect 166258 204892 166264 204904
rect 166316 204892 166322 204944
rect 65702 204280 65708 204332
rect 65760 204320 65766 204332
rect 68094 204320 68100 204332
rect 65760 204292 68100 204320
rect 65760 204280 65766 204292
rect 68094 204280 68100 204292
rect 68152 204280 68158 204332
rect 119798 204280 119804 204332
rect 119856 204320 119862 204332
rect 121454 204320 121460 204332
rect 119856 204292 121460 204320
rect 119856 204280 119862 204292
rect 121454 204280 121460 204292
rect 121512 204280 121518 204332
rect 233142 204280 233148 204332
rect 233200 204320 233206 204332
rect 580258 204320 580264 204332
rect 233200 204292 580264 204320
rect 233200 204280 233206 204292
rect 580258 204280 580264 204292
rect 580316 204280 580322 204332
rect 232682 204212 232688 204264
rect 232740 204252 232746 204264
rect 278038 204252 278044 204264
rect 232740 204224 278044 204252
rect 232740 204212 232746 204224
rect 278038 204212 278044 204224
rect 278096 204212 278102 204264
rect 126422 203532 126428 203584
rect 126480 203572 126486 203584
rect 167270 203572 167276 203584
rect 126480 203544 167276 203572
rect 126480 203532 126486 203544
rect 167270 203532 167276 203544
rect 167328 203532 167334 203584
rect 122558 202852 122564 202904
rect 122616 202892 122622 202904
rect 164970 202892 164976 202904
rect 122616 202864 164976 202892
rect 122616 202852 122622 202864
rect 164970 202852 164976 202864
rect 165028 202852 165034 202904
rect 232682 202784 232688 202836
rect 232740 202824 232746 202836
rect 289078 202824 289084 202836
rect 232740 202796 289084 202824
rect 232740 202784 232746 202796
rect 289078 202784 289084 202796
rect 289136 202784 289142 202836
rect 126330 202104 126336 202156
rect 126388 202144 126394 202156
rect 167454 202144 167460 202156
rect 126388 202116 167460 202144
rect 126388 202104 126394 202116
rect 167454 202104 167460 202116
rect 167512 202104 167518 202156
rect 3418 201492 3424 201544
rect 3476 201532 3482 201544
rect 63494 201532 63500 201544
rect 3476 201504 63500 201532
rect 3476 201492 3482 201504
rect 63494 201492 63500 201504
rect 63552 201492 63558 201544
rect 66714 201492 66720 201544
rect 66772 201532 66778 201544
rect 67634 201532 67640 201544
rect 66772 201504 67640 201532
rect 66772 201492 66778 201504
rect 67634 201492 67640 201504
rect 67692 201492 67698 201544
rect 121822 201492 121828 201544
rect 121880 201532 121886 201544
rect 124398 201532 124404 201544
rect 121880 201504 124404 201532
rect 121880 201492 121886 201504
rect 124398 201492 124404 201504
rect 124456 201492 124462 201544
rect 127710 201424 127716 201476
rect 127768 201464 127774 201476
rect 167086 201464 167092 201476
rect 127768 201436 167092 201464
rect 127768 201424 127774 201436
rect 167086 201424 167092 201436
rect 167144 201424 167150 201476
rect 167270 201152 167276 201204
rect 167328 201152 167334 201204
rect 167288 201000 167316 201152
rect 167270 200948 167276 201000
rect 167328 200948 167334 201000
rect 233326 200744 233332 200796
rect 233384 200784 233390 200796
rect 477494 200784 477500 200796
rect 233384 200756 477500 200784
rect 233384 200744 233390 200756
rect 477494 200744 477500 200756
rect 477552 200744 477558 200796
rect 119154 200512 119160 200524
rect 119080 200484 119160 200512
rect 69382 200336 69388 200388
rect 69440 200376 69446 200388
rect 72602 200376 72608 200388
rect 69440 200348 72608 200376
rect 69440 200336 69446 200348
rect 72602 200336 72608 200348
rect 72660 200336 72666 200388
rect 102824 200376 102830 200388
rect 98564 200348 102830 200376
rect 69842 200268 69848 200320
rect 69900 200308 69906 200320
rect 71268 200308 71274 200320
rect 69900 200280 71274 200308
rect 69900 200268 69906 200280
rect 71268 200268 71274 200280
rect 71326 200268 71332 200320
rect 73246 200268 73252 200320
rect 73304 200268 73310 200320
rect 74534 200268 74540 200320
rect 74592 200268 74598 200320
rect 75178 200308 75184 200320
rect 75104 200280 75184 200308
rect 67174 200132 67180 200184
rect 67232 200172 67238 200184
rect 69750 200172 69756 200184
rect 67232 200144 69756 200172
rect 67232 200132 67238 200144
rect 69750 200132 69756 200144
rect 69808 200132 69814 200184
rect 4798 200064 4804 200116
rect 4856 200104 4862 200116
rect 4856 200076 69704 200104
rect 4856 200064 4862 200076
rect 7558 199996 7564 200048
rect 7616 200036 7622 200048
rect 69566 200036 69572 200048
rect 7616 200008 69572 200036
rect 7616 199996 7622 200008
rect 69566 199996 69572 200008
rect 69624 199996 69630 200048
rect 69676 199968 69704 200076
rect 73264 199980 73292 200268
rect 74552 199980 74580 200268
rect 75104 199980 75132 200280
rect 75178 200268 75184 200280
rect 75236 200268 75242 200320
rect 76466 200268 76472 200320
rect 76524 200268 76530 200320
rect 77110 200268 77116 200320
rect 77168 200268 77174 200320
rect 77754 200268 77760 200320
rect 77812 200268 77818 200320
rect 79042 200268 79048 200320
rect 79100 200268 79106 200320
rect 79686 200268 79692 200320
rect 79744 200268 79750 200320
rect 80974 200268 80980 200320
rect 81032 200268 81038 200320
rect 81618 200268 81624 200320
rect 81676 200268 81682 200320
rect 82906 200268 82912 200320
rect 82964 200268 82970 200320
rect 83550 200268 83556 200320
rect 83608 200268 83614 200320
rect 84194 200268 84200 200320
rect 84252 200268 84258 200320
rect 85482 200268 85488 200320
rect 85540 200268 85546 200320
rect 86126 200268 86132 200320
rect 86184 200268 86190 200320
rect 87414 200268 87420 200320
rect 87472 200268 87478 200320
rect 88058 200308 88064 200320
rect 87984 200280 88064 200308
rect 76484 199980 76512 200268
rect 77128 199980 77156 200268
rect 77772 199980 77800 200268
rect 79060 199980 79088 200268
rect 79704 199980 79732 200268
rect 80992 199980 81020 200268
rect 81636 199980 81664 200268
rect 82924 199980 82952 200268
rect 83568 199980 83596 200268
rect 84212 199980 84240 200268
rect 85500 199980 85528 200268
rect 86144 199980 86172 200268
rect 87432 199980 87460 200268
rect 87984 199980 88012 200280
rect 88058 200268 88064 200280
rect 88116 200268 88122 200320
rect 89346 200268 89352 200320
rect 89404 200268 89410 200320
rect 89990 200268 89996 200320
rect 90048 200268 90054 200320
rect 90634 200268 90640 200320
rect 90692 200268 90698 200320
rect 91922 200308 91928 200320
rect 91848 200280 91928 200308
rect 89364 199980 89392 200268
rect 90008 200240 90036 200268
rect 89916 200212 90036 200240
rect 89916 199980 89944 200212
rect 90652 199980 90680 200268
rect 91848 199980 91876 200280
rect 91922 200268 91928 200280
rect 91980 200268 91986 200320
rect 92566 200268 92572 200320
rect 92624 200268 92630 200320
rect 93854 200268 93860 200320
rect 93912 200268 93918 200320
rect 94498 200308 94504 200320
rect 94424 200280 94504 200308
rect 92584 200240 92612 200268
rect 92492 200212 92612 200240
rect 92492 199980 92520 200212
rect 93872 199980 93900 200268
rect 94424 199980 94452 200280
rect 94498 200268 94504 200280
rect 94556 200268 94562 200320
rect 95786 200308 95792 200320
rect 95712 200280 95792 200308
rect 95712 199980 95740 200280
rect 95786 200268 95792 200280
rect 95844 200268 95850 200320
rect 96430 200268 96436 200320
rect 96488 200268 96494 200320
rect 97718 200268 97724 200320
rect 97776 200268 97782 200320
rect 98362 200308 98368 200320
rect 98288 200280 98368 200308
rect 96448 199980 96476 200268
rect 97736 200172 97764 200268
rect 97276 200144 97764 200172
rect 97276 199980 97304 200144
rect 98288 199980 98316 200280
rect 98362 200268 98368 200280
rect 98420 200268 98426 200320
rect 98564 199980 98592 200348
rect 102824 200336 102830 200348
rect 102882 200376 102888 200388
rect 102882 200348 104296 200376
rect 102882 200336 102888 200348
rect 99006 200268 99012 200320
rect 99064 200268 99070 200320
rect 100294 200268 100300 200320
rect 100352 200268 100358 200320
rect 100892 200268 100898 200320
rect 100950 200308 100956 200320
rect 100950 200280 101352 200308
rect 100950 200268 100956 200280
rect 99024 200172 99052 200268
rect 98932 200144 99052 200172
rect 98932 199980 98960 200144
rect 100312 199980 100340 200268
rect 101324 199980 101352 200280
rect 102226 200268 102232 200320
rect 102284 200268 102290 200320
rect 104158 200268 104164 200320
rect 104216 200268 104222 200320
rect 102244 200240 102272 200268
rect 102244 200212 102916 200240
rect 73154 199968 73160 199980
rect 69676 199940 73160 199968
rect 73154 199928 73160 199940
rect 73212 199928 73218 199980
rect 73246 199928 73252 199980
rect 73304 199928 73310 199980
rect 74534 199928 74540 199980
rect 74592 199928 74598 199980
rect 75086 199928 75092 199980
rect 75144 199928 75150 199980
rect 76466 199928 76472 199980
rect 76524 199928 76530 199980
rect 77110 199928 77116 199980
rect 77168 199928 77174 199980
rect 77754 199928 77760 199980
rect 77812 199928 77818 199980
rect 79042 199928 79048 199980
rect 79100 199928 79106 199980
rect 79686 199928 79692 199980
rect 79744 199928 79750 199980
rect 80974 199928 80980 199980
rect 81032 199928 81038 199980
rect 81618 199928 81624 199980
rect 81676 199928 81682 199980
rect 82906 199928 82912 199980
rect 82964 199928 82970 199980
rect 83550 199928 83556 199980
rect 83608 199928 83614 199980
rect 84194 199928 84200 199980
rect 84252 199928 84258 199980
rect 85482 199928 85488 199980
rect 85540 199928 85546 199980
rect 86126 199928 86132 199980
rect 86184 199928 86190 199980
rect 87414 199928 87420 199980
rect 87472 199928 87478 199980
rect 87966 199928 87972 199980
rect 88024 199928 88030 199980
rect 89346 199928 89352 199980
rect 89404 199928 89410 199980
rect 89898 199928 89904 199980
rect 89956 199928 89962 199980
rect 90634 199928 90640 199980
rect 90692 199928 90698 199980
rect 91830 199928 91836 199980
rect 91888 199928 91894 199980
rect 92474 199928 92480 199980
rect 92532 199928 92538 199980
rect 93854 199928 93860 199980
rect 93912 199928 93918 199980
rect 94406 199928 94412 199980
rect 94464 199928 94470 199980
rect 95694 199928 95700 199980
rect 95752 199928 95758 199980
rect 96430 199928 96436 199980
rect 96488 199928 96494 199980
rect 97258 199928 97264 199980
rect 97316 199928 97322 199980
rect 98270 199928 98276 199980
rect 98328 199928 98334 199980
rect 98546 199928 98552 199980
rect 98604 199928 98610 199980
rect 98914 199928 98920 199980
rect 98972 199928 98978 199980
rect 100294 199928 100300 199980
rect 100352 199928 100358 199980
rect 101306 199928 101312 199980
rect 101364 199928 101370 199980
rect 102888 199968 102916 200212
rect 104176 199980 104204 200268
rect 104268 199980 104296 200348
rect 111242 200336 111248 200388
rect 111300 200376 111306 200388
rect 111300 200348 111380 200376
rect 111300 200336 111306 200348
rect 104802 200268 104808 200320
rect 104860 200268 104866 200320
rect 105400 200268 105406 200320
rect 105458 200268 105464 200320
rect 106734 200268 106740 200320
rect 106792 200268 106798 200320
rect 107378 200268 107384 200320
rect 107436 200308 107442 200320
rect 107436 200280 107516 200308
rect 107436 200268 107442 200280
rect 104820 199980 104848 200268
rect 105418 199980 105446 200268
rect 106752 200104 106780 200268
rect 103422 199968 103428 199980
rect 102888 199940 103428 199968
rect 103422 199928 103428 199940
rect 103480 199928 103486 199980
rect 104158 199928 104164 199980
rect 104216 199928 104222 199980
rect 104250 199928 104256 199980
rect 104308 199928 104314 199980
rect 104802 199928 104808 199980
rect 104860 199928 104866 199980
rect 105354 199928 105360 199980
rect 105412 199940 105446 199980
rect 106476 200076 106780 200104
rect 105412 199928 105418 199940
rect 64506 199860 64512 199912
rect 64564 199900 64570 199912
rect 75178 199900 75184 199912
rect 64564 199872 75184 199900
rect 64564 199860 64570 199872
rect 75178 199860 75184 199872
rect 75236 199860 75242 199912
rect 84654 199860 84660 199912
rect 84712 199900 84718 199912
rect 101324 199900 101352 199928
rect 84712 199872 101352 199900
rect 84712 199860 84718 199872
rect 62758 199792 62764 199844
rect 62816 199832 62822 199844
rect 62816 199804 80054 199832
rect 62816 199792 62822 199804
rect 61378 199724 61384 199776
rect 61436 199764 61442 199776
rect 75270 199764 75276 199776
rect 61436 199736 75276 199764
rect 61436 199724 61442 199736
rect 75270 199724 75276 199736
rect 75328 199724 75334 199776
rect 80026 199764 80054 199804
rect 84838 199792 84844 199844
rect 84896 199832 84902 199844
rect 98638 199832 98644 199844
rect 84896 199804 98644 199832
rect 84896 199792 84902 199804
rect 98638 199792 98644 199804
rect 98696 199792 98702 199844
rect 106476 199832 106504 200076
rect 107488 199980 107516 200280
rect 108666 200268 108672 200320
rect 108724 200268 108730 200320
rect 109310 200268 109316 200320
rect 109368 200268 109374 200320
rect 110598 200268 110604 200320
rect 110656 200308 110662 200320
rect 110656 200280 111288 200308
rect 110656 200268 110662 200280
rect 107470 199928 107476 199980
rect 107528 199928 107534 199980
rect 108684 199968 108712 200268
rect 109328 199980 109356 200268
rect 111260 199980 111288 200280
rect 108758 199968 108764 199980
rect 108684 199940 108764 199968
rect 108758 199928 108764 199940
rect 108816 199928 108822 199980
rect 109310 199928 109316 199980
rect 109368 199928 109374 199980
rect 111242 199928 111248 199980
rect 111300 199928 111306 199980
rect 111150 199860 111156 199912
rect 111208 199900 111214 199912
rect 111352 199900 111380 200348
rect 113174 200336 113180 200388
rect 113232 200376 113238 200388
rect 113232 200348 114508 200376
rect 113232 200336 113238 200348
rect 111886 200268 111892 200320
rect 111944 200268 111950 200320
rect 113772 200308 113778 200320
rect 113192 200280 113778 200308
rect 111904 200104 111932 200268
rect 111904 200076 112576 200104
rect 112548 199980 112576 200076
rect 113192 199980 113220 200280
rect 113772 200268 113778 200280
rect 113830 200268 113836 200320
rect 114480 199980 114508 200348
rect 115106 200268 115112 200320
rect 115164 200308 115170 200320
rect 115164 200280 115336 200308
rect 115164 200268 115170 200280
rect 115308 199980 115336 200280
rect 115750 200268 115756 200320
rect 115808 200308 115814 200320
rect 115808 200280 115888 200308
rect 115808 200268 115814 200280
rect 115860 199980 115888 200280
rect 117038 200268 117044 200320
rect 117096 200268 117102 200320
rect 117682 200268 117688 200320
rect 117740 200268 117746 200320
rect 112530 199928 112536 199980
rect 112588 199928 112594 199980
rect 113174 199928 113180 199980
rect 113232 199928 113238 199980
rect 114462 199928 114468 199980
rect 114520 199928 114526 199980
rect 115290 199928 115296 199980
rect 115348 199928 115354 199980
rect 115842 199928 115848 199980
rect 115900 199928 115906 199980
rect 116578 199928 116584 199980
rect 116636 199968 116642 199980
rect 117056 199968 117084 200268
rect 117700 200036 117728 200268
rect 119080 200116 119108 200484
rect 119154 200472 119160 200484
rect 119212 200472 119218 200524
rect 122558 200132 122564 200184
rect 122616 200172 122622 200184
rect 152550 200172 152556 200184
rect 122616 200144 152556 200172
rect 122616 200132 122622 200144
rect 152550 200132 152556 200144
rect 152608 200132 152614 200184
rect 119062 200064 119068 200116
rect 119120 200064 119126 200116
rect 117332 200008 117728 200036
rect 117332 199980 117360 200008
rect 116636 199940 117084 199968
rect 116636 199928 116642 199940
rect 117314 199928 117320 199980
rect 117372 199928 117378 199980
rect 117682 199928 117688 199980
rect 117740 199968 117746 199980
rect 138014 199968 138020 199980
rect 117740 199940 138020 199968
rect 117740 199928 117746 199940
rect 138014 199928 138020 199940
rect 138072 199928 138078 199980
rect 111208 199872 111380 199900
rect 111208 199860 111214 199872
rect 107194 199832 107200 199844
rect 99346 199804 107200 199832
rect 98730 199764 98736 199776
rect 80026 199736 98736 199764
rect 98730 199724 98736 199736
rect 98788 199724 98794 199776
rect 65518 199656 65524 199708
rect 65576 199696 65582 199708
rect 74810 199696 74816 199708
rect 65576 199668 74816 199696
rect 65576 199656 65582 199668
rect 74810 199656 74816 199668
rect 74868 199656 74874 199708
rect 74994 199656 75000 199708
rect 75052 199696 75058 199708
rect 99346 199696 99374 199804
rect 107194 199792 107200 199804
rect 107252 199792 107258 199844
rect 112530 199764 112536 199776
rect 75052 199668 99374 199696
rect 104176 199736 112536 199764
rect 75052 199656 75058 199668
rect 69566 199588 69572 199640
rect 69624 199628 69630 199640
rect 74718 199628 74724 199640
rect 69624 199600 74724 199628
rect 69624 199588 69630 199600
rect 74718 199588 74724 199600
rect 74776 199588 74782 199640
rect 75270 199588 75276 199640
rect 75328 199628 75334 199640
rect 104176 199628 104204 199736
rect 112530 199724 112536 199736
rect 112588 199724 112594 199776
rect 113818 199724 113824 199776
rect 113876 199764 113882 199776
rect 125042 199764 125048 199776
rect 113876 199736 125048 199764
rect 113876 199724 113882 199736
rect 125042 199724 125048 199736
rect 125100 199724 125106 199776
rect 108114 199656 108120 199708
rect 108172 199696 108178 199708
rect 120074 199696 120080 199708
rect 108172 199668 120080 199696
rect 108172 199656 108178 199668
rect 120074 199656 120080 199668
rect 120132 199656 120138 199708
rect 75328 199600 104204 199628
rect 75328 199588 75334 199600
rect 108666 199588 108672 199640
rect 108724 199628 108730 199640
rect 120442 199628 120448 199640
rect 108724 199600 120448 199628
rect 108724 199588 108730 199600
rect 120442 199588 120448 199600
rect 120500 199588 120506 199640
rect 68738 199520 68744 199572
rect 68796 199560 68802 199572
rect 157334 199560 157340 199572
rect 68796 199532 157340 199560
rect 68796 199520 68802 199532
rect 157334 199520 157340 199532
rect 157392 199520 157398 199572
rect 69014 199452 69020 199504
rect 69072 199492 69078 199504
rect 167362 199492 167368 199504
rect 69072 199464 167368 199492
rect 69072 199452 69078 199464
rect 167362 199452 167368 199464
rect 167420 199452 167426 199504
rect 65610 199384 65616 199436
rect 65668 199424 65674 199436
rect 168190 199424 168196 199436
rect 65668 199396 168196 199424
rect 65668 199384 65674 199396
rect 168190 199384 168196 199396
rect 168248 199424 168254 199436
rect 169018 199424 169024 199436
rect 168248 199396 169024 199424
rect 168248 199384 168254 199396
rect 169018 199384 169024 199396
rect 169076 199384 169082 199436
rect 67910 199316 67916 199368
rect 67968 199356 67974 199368
rect 72694 199356 72700 199368
rect 67968 199328 72700 199356
rect 67968 199316 67974 199328
rect 72694 199316 72700 199328
rect 72752 199316 72758 199368
rect 73154 199316 73160 199368
rect 73212 199356 73218 199368
rect 84746 199356 84752 199368
rect 73212 199328 84752 199356
rect 73212 199316 73218 199328
rect 84746 199316 84752 199328
rect 84804 199316 84810 199368
rect 84930 199316 84936 199368
rect 84988 199356 84994 199368
rect 84988 199328 98684 199356
rect 84988 199316 84994 199328
rect 75178 199248 75184 199300
rect 75236 199288 75242 199300
rect 82078 199288 82084 199300
rect 75236 199260 82084 199288
rect 75236 199248 75242 199260
rect 82078 199248 82084 199260
rect 82136 199248 82142 199300
rect 98546 199288 98552 199300
rect 89686 199260 98552 199288
rect 74718 199180 74724 199232
rect 74776 199220 74782 199232
rect 84654 199220 84660 199232
rect 74776 199192 84660 199220
rect 74776 199180 74782 199192
rect 84654 199180 84660 199192
rect 84712 199180 84718 199232
rect 84746 199180 84752 199232
rect 84804 199220 84810 199232
rect 89686 199220 89714 199260
rect 98546 199248 98552 199260
rect 98604 199248 98610 199300
rect 98656 199288 98684 199328
rect 98730 199316 98736 199368
rect 98788 199356 98794 199368
rect 113726 199356 113732 199368
rect 98788 199328 113732 199356
rect 98788 199316 98794 199328
rect 113726 199316 113732 199328
rect 113784 199316 113790 199368
rect 113818 199288 113824 199300
rect 98656 199260 113824 199288
rect 113818 199248 113824 199260
rect 113876 199248 113882 199300
rect 84804 199192 89714 199220
rect 84804 199180 84810 199192
rect 98638 199180 98644 199232
rect 98696 199220 98702 199232
rect 117682 199220 117688 199232
rect 98696 199192 117688 199220
rect 98696 199180 98702 199192
rect 117682 199180 117688 199192
rect 117740 199180 117746 199232
rect 65794 199112 65800 199164
rect 65852 199152 65858 199164
rect 84838 199152 84844 199164
rect 65852 199124 84844 199152
rect 65852 199112 65858 199124
rect 84838 199112 84844 199124
rect 84896 199112 84902 199164
rect 117130 198908 117136 198960
rect 117188 198948 117194 198960
rect 122374 198948 122380 198960
rect 117188 198920 122380 198948
rect 117188 198908 117194 198920
rect 122374 198908 122380 198920
rect 122432 198908 122438 198960
rect 117222 198840 117228 198892
rect 117280 198880 117286 198892
rect 122006 198880 122012 198892
rect 117280 198852 122012 198880
rect 117280 198840 117286 198852
rect 122006 198840 122012 198852
rect 122064 198840 122070 198892
rect 117038 198772 117044 198824
rect 117096 198812 117102 198824
rect 121638 198812 121644 198824
rect 117096 198784 121644 198812
rect 117096 198772 117102 198784
rect 121638 198772 121644 198784
rect 121696 198772 121702 198824
rect 68830 198704 68836 198756
rect 68888 198744 68894 198756
rect 71038 198744 71044 198756
rect 68888 198716 71044 198744
rect 68888 198704 68894 198716
rect 71038 198704 71044 198716
rect 71096 198704 71102 198756
rect 118510 198704 118516 198756
rect 118568 198744 118574 198756
rect 121546 198744 121552 198756
rect 118568 198716 121552 198744
rect 118568 198704 118574 198716
rect 121546 198704 121552 198716
rect 121604 198704 121610 198756
rect 68554 198636 68560 198688
rect 68612 198676 68618 198688
rect 164878 198676 164884 198688
rect 68612 198648 164884 198676
rect 68612 198636 68618 198648
rect 164878 198636 164884 198648
rect 164936 198636 164942 198688
rect 18598 198568 18604 198620
rect 18656 198608 18662 198620
rect 87414 198608 87420 198620
rect 18656 198580 87420 198608
rect 18656 198568 18662 198580
rect 87414 198568 87420 198580
rect 87472 198568 87478 198620
rect 91830 198568 91836 198620
rect 91888 198608 91894 198620
rect 91888 198580 104204 198608
rect 91888 198568 91894 198580
rect 58618 198500 58624 198552
rect 58676 198540 58682 198552
rect 104066 198540 104072 198552
rect 58676 198512 104072 198540
rect 58676 198500 58682 198512
rect 104066 198500 104072 198512
rect 104124 198500 104130 198552
rect 104176 198540 104204 198580
rect 108758 198568 108764 198620
rect 108816 198608 108822 198620
rect 110414 198608 110420 198620
rect 108816 198580 110420 198608
rect 108816 198568 108822 198580
rect 110414 198568 110420 198580
rect 110472 198568 110478 198620
rect 104176 198512 109034 198540
rect 55858 198432 55864 198484
rect 55916 198472 55922 198484
rect 97258 198472 97264 198484
rect 55916 198444 97264 198472
rect 55916 198432 55922 198444
rect 97258 198432 97264 198444
rect 97316 198432 97322 198484
rect 98914 198432 98920 198484
rect 98972 198472 98978 198484
rect 106274 198472 106280 198484
rect 98972 198444 106280 198472
rect 98972 198432 98978 198444
rect 106274 198432 106280 198444
rect 106332 198432 106338 198484
rect 109006 198472 109034 198512
rect 113818 198500 113824 198552
rect 113876 198540 113882 198552
rect 117314 198540 117320 198552
rect 113876 198512 117320 198540
rect 113876 198500 113882 198512
rect 117314 198500 117320 198512
rect 117372 198500 117378 198552
rect 111794 198472 111800 198484
rect 109006 198444 111800 198472
rect 111794 198432 111800 198444
rect 111852 198432 111858 198484
rect 66162 198364 66168 198416
rect 66220 198404 66226 198416
rect 75086 198404 75092 198416
rect 66220 198376 75092 198404
rect 66220 198364 66226 198376
rect 75086 198364 75092 198376
rect 75144 198364 75150 198416
rect 81618 198364 81624 198416
rect 81676 198404 81682 198416
rect 106918 198404 106924 198416
rect 81676 198376 106924 198404
rect 81676 198364 81682 198376
rect 106918 198364 106924 198376
rect 106976 198364 106982 198416
rect 107194 198364 107200 198416
rect 107252 198404 107258 198416
rect 127066 198404 127072 198416
rect 107252 198376 127072 198404
rect 107252 198364 107258 198376
rect 127066 198364 127072 198376
rect 127124 198364 127130 198416
rect 101306 198296 101312 198348
rect 101364 198336 101370 198348
rect 129734 198336 129740 198348
rect 101364 198308 129740 198336
rect 101364 198296 101370 198308
rect 129734 198296 129740 198308
rect 129792 198296 129798 198348
rect 104250 198228 104256 198280
rect 104308 198268 104314 198280
rect 131114 198268 131120 198280
rect 104308 198240 131120 198268
rect 104308 198228 104314 198240
rect 131114 198228 131120 198240
rect 131172 198228 131178 198280
rect 65794 198160 65800 198212
rect 65852 198200 65858 198212
rect 79042 198200 79048 198212
rect 65852 198172 79048 198200
rect 65852 198160 65858 198172
rect 79042 198160 79048 198172
rect 79100 198160 79106 198212
rect 95694 198160 95700 198212
rect 95752 198200 95758 198212
rect 126330 198200 126336 198212
rect 95752 198172 126336 198200
rect 95752 198160 95758 198172
rect 126330 198160 126336 198172
rect 126388 198160 126394 198212
rect 63218 198092 63224 198144
rect 63276 198132 63282 198144
rect 69382 198132 69388 198144
rect 63276 198104 69388 198132
rect 63276 198092 63282 198104
rect 69382 198092 69388 198104
rect 69440 198092 69446 198144
rect 107470 198092 107476 198144
rect 107528 198132 107534 198144
rect 137278 198132 137284 198144
rect 107528 198104 137284 198132
rect 107528 198092 107534 198104
rect 137278 198092 137284 198104
rect 137336 198092 137342 198144
rect 157334 198092 157340 198144
rect 157392 198132 157398 198144
rect 158162 198132 158168 198144
rect 157392 198104 158168 198132
rect 157392 198092 157398 198104
rect 158162 198092 158168 198104
rect 158220 198132 158226 198144
rect 167362 198132 167368 198144
rect 158220 198104 167368 198132
rect 158220 198092 158226 198104
rect 167362 198092 167368 198104
rect 167420 198092 167426 198144
rect 61838 198024 61844 198076
rect 61896 198064 61902 198076
rect 79686 198064 79692 198076
rect 61896 198036 79692 198064
rect 61896 198024 61902 198036
rect 79686 198024 79692 198036
rect 79744 198024 79750 198076
rect 85482 198024 85488 198076
rect 85540 198064 85546 198076
rect 111058 198064 111064 198076
rect 85540 198036 111064 198064
rect 85540 198024 85546 198036
rect 111058 198024 111064 198036
rect 111116 198024 111122 198076
rect 114462 198024 114468 198076
rect 114520 198064 114526 198076
rect 170306 198064 170312 198076
rect 114520 198036 170312 198064
rect 114520 198024 114526 198036
rect 170306 198024 170312 198036
rect 170364 198024 170370 198076
rect 65886 197956 65892 198008
rect 65944 197996 65950 198008
rect 168282 197996 168288 198008
rect 65944 197968 168288 197996
rect 65944 197956 65950 197968
rect 168282 197956 168288 197968
rect 168340 197996 168346 198008
rect 169754 197996 169760 198008
rect 168340 197968 169760 197996
rect 168340 197956 168346 197968
rect 169754 197956 169760 197968
rect 169812 197956 169818 198008
rect 86126 197888 86132 197940
rect 86184 197928 86190 197940
rect 109034 197928 109040 197940
rect 86184 197900 109040 197928
rect 86184 197888 86190 197900
rect 109034 197888 109040 197900
rect 109092 197888 109098 197940
rect 77110 197820 77116 197872
rect 77168 197860 77174 197872
rect 79318 197860 79324 197872
rect 77168 197832 79324 197860
rect 77168 197820 77174 197832
rect 79318 197820 79324 197832
rect 79376 197820 79382 197872
rect 89898 197820 89904 197872
rect 89956 197860 89962 197872
rect 108390 197860 108396 197872
rect 89956 197832 108396 197860
rect 89956 197820 89962 197832
rect 108390 197820 108396 197832
rect 108448 197820 108454 197872
rect 104066 197752 104072 197804
rect 104124 197792 104130 197804
rect 111150 197792 111156 197804
rect 104124 197764 111156 197792
rect 104124 197752 104130 197764
rect 111150 197752 111156 197764
rect 111208 197752 111214 197804
rect 104802 197684 104808 197736
rect 104860 197724 104866 197736
rect 109126 197724 109132 197736
rect 104860 197696 109132 197724
rect 104860 197684 104866 197696
rect 109126 197684 109132 197696
rect 109184 197684 109190 197736
rect 104158 197616 104164 197668
rect 104216 197656 104222 197668
rect 110506 197656 110512 197668
rect 104216 197628 110512 197656
rect 104216 197616 104222 197628
rect 110506 197616 110512 197628
rect 110564 197616 110570 197668
rect 137278 197616 137284 197668
rect 137336 197656 137342 197668
rect 166350 197656 166356 197668
rect 137336 197628 166356 197656
rect 137336 197616 137342 197628
rect 166350 197616 166356 197628
rect 166408 197616 166414 197668
rect 131114 197548 131120 197600
rect 131172 197588 131178 197600
rect 131758 197588 131764 197600
rect 131172 197560 131764 197588
rect 131172 197548 131178 197560
rect 131758 197548 131764 197560
rect 131816 197588 131822 197600
rect 166442 197588 166448 197600
rect 131816 197560 166448 197588
rect 131816 197548 131822 197560
rect 166442 197548 166448 197560
rect 166500 197548 166506 197600
rect 126330 197480 126336 197532
rect 126388 197520 126394 197532
rect 166258 197520 166264 197532
rect 126388 197492 166264 197520
rect 126388 197480 126394 197492
rect 166258 197480 166264 197492
rect 166316 197480 166322 197532
rect 117958 197412 117964 197464
rect 118016 197452 118022 197464
rect 119154 197452 119160 197464
rect 118016 197424 119160 197452
rect 118016 197412 118022 197424
rect 119154 197412 119160 197424
rect 119212 197412 119218 197464
rect 129734 197412 129740 197464
rect 129792 197452 129798 197464
rect 130378 197452 130384 197464
rect 129792 197424 130384 197452
rect 129792 197412 129798 197424
rect 130378 197412 130384 197424
rect 130436 197452 130442 197464
rect 170398 197452 170404 197464
rect 130436 197424 170404 197452
rect 130436 197412 130442 197424
rect 170398 197412 170404 197424
rect 170456 197412 170462 197464
rect 92474 197344 92480 197396
rect 92532 197384 92538 197396
rect 94590 197384 94596 197396
rect 92532 197356 94596 197384
rect 92532 197344 92538 197356
rect 94590 197344 94596 197356
rect 94648 197344 94654 197396
rect 118602 197344 118608 197396
rect 118660 197384 118666 197396
rect 119614 197384 119620 197396
rect 118660 197356 119620 197384
rect 118660 197344 118666 197356
rect 119614 197344 119620 197356
rect 119672 197344 119678 197396
rect 127066 197344 127072 197396
rect 127124 197384 127130 197396
rect 127710 197384 127716 197396
rect 127124 197356 127716 197384
rect 127124 197344 127130 197356
rect 127710 197344 127716 197356
rect 127768 197384 127774 197396
rect 170490 197384 170496 197396
rect 127768 197356 170496 197384
rect 127768 197344 127774 197356
rect 170490 197344 170496 197356
rect 170548 197344 170554 197396
rect 76466 196732 76472 196784
rect 76524 196772 76530 196784
rect 86218 196772 86224 196784
rect 76524 196744 86224 196772
rect 76524 196732 76530 196744
rect 86218 196732 86224 196744
rect 86276 196732 86282 196784
rect 108758 196732 108764 196784
rect 108816 196772 108822 196784
rect 119430 196772 119436 196784
rect 108816 196744 119436 196772
rect 108816 196732 108822 196744
rect 119430 196732 119436 196744
rect 119488 196732 119494 196784
rect 69106 196664 69112 196716
rect 69164 196704 69170 196716
rect 128354 196704 128360 196716
rect 69164 196676 128360 196704
rect 69164 196664 69170 196676
rect 128354 196664 128360 196676
rect 128412 196664 128418 196716
rect 69474 196596 69480 196648
rect 69532 196636 69538 196648
rect 70302 196636 70308 196648
rect 69532 196608 70308 196636
rect 69532 196596 69538 196608
rect 70302 196596 70308 196608
rect 70360 196636 70366 196648
rect 167362 196636 167368 196648
rect 70360 196608 167368 196636
rect 70360 196596 70366 196608
rect 167362 196596 167368 196608
rect 167420 196596 167426 196648
rect 118694 195984 118700 196036
rect 118752 196024 118758 196036
rect 119706 196024 119712 196036
rect 118752 195996 119712 196024
rect 118752 195984 118758 195996
rect 119706 195984 119712 195996
rect 119764 196024 119770 196036
rect 169018 196024 169024 196036
rect 119764 195996 169024 196024
rect 119764 195984 119770 195996
rect 169018 195984 169024 195996
rect 169076 195984 169082 196036
rect 105354 195508 105360 195560
rect 105412 195548 105418 195560
rect 113266 195548 113272 195560
rect 105412 195520 113272 195548
rect 105412 195508 105418 195520
rect 113266 195508 113272 195520
rect 113324 195508 113330 195560
rect 100294 195440 100300 195492
rect 100352 195480 100358 195492
rect 110598 195480 110604 195492
rect 100352 195452 110604 195480
rect 100352 195440 100358 195452
rect 110598 195440 110604 195452
rect 110656 195440 110662 195492
rect 98270 195372 98276 195424
rect 98328 195412 98334 195424
rect 113358 195412 113364 195424
rect 98328 195384 113364 195412
rect 98328 195372 98334 195384
rect 113358 195372 113364 195384
rect 113416 195372 113422 195424
rect 94406 195304 94412 195356
rect 94464 195344 94470 195356
rect 115934 195344 115940 195356
rect 94464 195316 115940 195344
rect 94464 195304 94470 195316
rect 115934 195304 115940 195316
rect 115992 195304 115998 195356
rect 87966 195236 87972 195288
rect 88024 195276 88030 195288
rect 114554 195276 114560 195288
rect 88024 195248 114560 195276
rect 88024 195236 88030 195248
rect 114554 195236 114560 195248
rect 114612 195236 114618 195288
rect 115658 194896 115664 194948
rect 115716 194936 115722 194948
rect 121914 194936 121920 194948
rect 115716 194908 121920 194936
rect 115716 194896 115722 194908
rect 121914 194896 121920 194908
rect 121972 194896 121978 194948
rect 116578 194624 116584 194676
rect 116636 194664 116642 194676
rect 166534 194664 166540 194676
rect 116636 194636 166540 194664
rect 116636 194624 116642 194636
rect 166534 194624 166540 194636
rect 166592 194624 166598 194676
rect 3418 194556 3424 194608
rect 3476 194596 3482 194608
rect 117958 194596 117964 194608
rect 3476 194568 117964 194596
rect 3476 194556 3482 194568
rect 117958 194556 117964 194568
rect 118016 194556 118022 194608
rect 113082 193944 113088 193996
rect 113140 193984 113146 193996
rect 118694 193984 118700 193996
rect 113140 193956 118700 193984
rect 113140 193944 113146 193956
rect 118694 193944 118700 193956
rect 118752 193944 118758 193996
rect 108482 193876 108488 193928
rect 108540 193916 108546 193928
rect 120166 193916 120172 193928
rect 108540 193888 120172 193916
rect 108540 193876 108546 193888
rect 120166 193876 120172 193888
rect 120224 193876 120230 193928
rect 63494 193808 63500 193860
rect 63552 193848 63558 193860
rect 111886 193848 111892 193860
rect 63552 193820 111892 193848
rect 63552 193808 63558 193820
rect 111886 193808 111892 193820
rect 111944 193848 111950 193860
rect 122098 193848 122104 193860
rect 111944 193820 122104 193848
rect 111944 193808 111950 193820
rect 122098 193808 122104 193820
rect 122156 193808 122162 193860
rect 115750 193672 115756 193724
rect 115808 193712 115814 193724
rect 122742 193712 122748 193724
rect 115808 193684 122748 193712
rect 115808 193672 115814 193684
rect 122742 193672 122748 193684
rect 122800 193672 122806 193724
rect 68462 192448 68468 192500
rect 68520 192488 68526 192500
rect 167362 192488 167368 192500
rect 68520 192460 167368 192488
rect 68520 192448 68526 192460
rect 167362 192448 167368 192460
rect 167420 192448 167426 192500
rect 233878 191836 233884 191888
rect 233936 191876 233942 191888
rect 579706 191876 579712 191888
rect 233936 191848 579712 191876
rect 233936 191836 233942 191848
rect 579706 191836 579712 191848
rect 579764 191836 579770 191888
rect 66806 191088 66812 191140
rect 66864 191128 66870 191140
rect 168098 191128 168104 191140
rect 66864 191100 168104 191128
rect 66864 191088 66870 191100
rect 168098 191088 168104 191100
rect 168156 191088 168162 191140
rect 233142 191088 233148 191140
rect 233200 191128 233206 191140
rect 233418 191128 233424 191140
rect 233200 191100 233424 191128
rect 233200 191088 233206 191100
rect 233418 191088 233424 191100
rect 233476 191128 233482 191140
rect 578878 191128 578884 191140
rect 233476 191100 578884 191128
rect 233476 191088 233482 191100
rect 578878 191088 578884 191100
rect 578936 191088 578942 191140
rect 115842 190544 115848 190596
rect 115900 190584 115906 190596
rect 115900 190556 122834 190584
rect 115900 190544 115906 190556
rect 113818 190476 113824 190528
rect 113876 190516 113882 190528
rect 118050 190516 118056 190528
rect 113876 190488 118056 190516
rect 113876 190476 113882 190488
rect 118050 190476 118056 190488
rect 118108 190476 118114 190528
rect 122806 190516 122834 190556
rect 162394 190516 162400 190528
rect 122806 190488 162400 190516
rect 162394 190476 162400 190488
rect 162452 190476 162458 190528
rect 89346 189796 89352 189848
rect 89404 189836 89410 189848
rect 123478 189836 123484 189848
rect 89404 189808 123484 189836
rect 89404 189796 89410 189808
rect 123478 189796 123484 189808
rect 123536 189796 123542 189848
rect 64414 189728 64420 189780
rect 64472 189768 64478 189780
rect 155862 189768 155868 189780
rect 64472 189740 155868 189768
rect 64472 189728 64478 189740
rect 155862 189728 155868 189740
rect 155920 189728 155926 189780
rect 142982 189116 142988 189168
rect 143040 189156 143046 189168
rect 144270 189156 144276 189168
rect 143040 189128 144276 189156
rect 143040 189116 143046 189128
rect 144270 189116 144276 189128
rect 144328 189116 144334 189168
rect 155862 189116 155868 189168
rect 155920 189156 155926 189168
rect 167362 189156 167368 189168
rect 155920 189128 167368 189156
rect 155920 189116 155926 189128
rect 167362 189116 167368 189128
rect 167420 189116 167426 189168
rect 123478 189048 123484 189100
rect 123536 189088 123542 189100
rect 164878 189088 164884 189100
rect 123536 189060 164884 189088
rect 123536 189048 123542 189060
rect 164878 189048 164884 189060
rect 164936 189048 164942 189100
rect 110230 188300 110236 188352
rect 110288 188340 110294 188352
rect 122650 188340 122656 188352
rect 110288 188312 122656 188340
rect 110288 188300 110294 188312
rect 122650 188300 122656 188312
rect 122708 188300 122714 188352
rect 233142 188300 233148 188352
rect 233200 188340 233206 188352
rect 233510 188340 233516 188352
rect 233200 188312 233516 188340
rect 233200 188300 233206 188312
rect 233510 188300 233516 188312
rect 233568 188340 233574 188352
rect 242158 188340 242164 188352
rect 233568 188312 242164 188340
rect 233568 188300 233574 188312
rect 242158 188300 242164 188312
rect 242216 188300 242222 188352
rect 72694 186940 72700 186992
rect 72752 186980 72758 186992
rect 150526 186980 150532 186992
rect 72752 186952 150532 186980
rect 72752 186940 72758 186952
rect 150526 186940 150532 186952
rect 150584 186940 150590 186992
rect 233142 186940 233148 186992
rect 233200 186980 233206 186992
rect 233602 186980 233608 186992
rect 233200 186952 233608 186980
rect 233200 186940 233206 186952
rect 233602 186940 233608 186952
rect 233660 186980 233666 186992
rect 249058 186980 249064 186992
rect 233660 186952 249064 186980
rect 233660 186940 233666 186952
rect 249058 186940 249064 186952
rect 249116 186940 249122 186992
rect 150526 186328 150532 186380
rect 150584 186368 150590 186380
rect 151722 186368 151728 186380
rect 150584 186340 151728 186368
rect 150584 186328 150590 186340
rect 151722 186328 151728 186340
rect 151780 186368 151786 186380
rect 167362 186368 167368 186380
rect 151780 186340 167368 186368
rect 151780 186328 151786 186340
rect 167362 186328 167368 186340
rect 167420 186328 167426 186380
rect 69658 185580 69664 185632
rect 69716 185620 69722 185632
rect 167362 185620 167368 185632
rect 69716 185592 167368 185620
rect 69716 185580 69722 185592
rect 167362 185580 167368 185592
rect 167420 185580 167426 185632
rect 68002 184832 68008 184884
rect 68060 184872 68066 184884
rect 167362 184872 167368 184884
rect 68060 184844 167368 184872
rect 68060 184832 68066 184844
rect 167362 184832 167368 184844
rect 167420 184832 167426 184884
rect 82906 184152 82912 184204
rect 82964 184192 82970 184204
rect 116670 184192 116676 184204
rect 82964 184164 116676 184192
rect 82964 184152 82970 184164
rect 116670 184152 116676 184164
rect 116728 184152 116734 184204
rect 116670 183540 116676 183592
rect 116728 183580 116734 183592
rect 156874 183580 156880 183592
rect 116728 183552 156880 183580
rect 116728 183540 116734 183552
rect 156874 183540 156880 183552
rect 156932 183540 156938 183592
rect 72602 183472 72608 183524
rect 72660 183512 72666 183524
rect 167362 183512 167368 183524
rect 72660 183484 167368 183512
rect 72660 183472 72666 183484
rect 167362 183472 167368 183484
rect 167420 183472 167426 183524
rect 110322 183404 110328 183456
rect 110380 183444 110386 183456
rect 115290 183444 115296 183456
rect 110380 183416 115296 183444
rect 110380 183404 110386 183416
rect 115290 183404 115296 183416
rect 115348 183404 115354 183456
rect 117958 183404 117964 183456
rect 118016 183444 118022 183456
rect 123846 183444 123852 183456
rect 118016 183416 123852 183444
rect 118016 183404 118022 183416
rect 123846 183404 123852 183416
rect 123904 183404 123910 183456
rect 90634 182792 90640 182844
rect 90692 182832 90698 182844
rect 123478 182832 123484 182844
rect 90692 182804 123484 182832
rect 90692 182792 90698 182804
rect 123478 182792 123484 182804
rect 123536 182792 123542 182844
rect 123478 182180 123484 182232
rect 123536 182220 123542 182232
rect 163498 182220 163504 182232
rect 123536 182192 163504 182220
rect 123536 182180 123542 182192
rect 163498 182180 163504 182192
rect 163556 182180 163562 182232
rect 77754 181432 77760 181484
rect 77812 181472 77818 181484
rect 112438 181472 112444 181484
rect 77812 181444 112444 181472
rect 77812 181432 77818 181444
rect 112438 181432 112444 181444
rect 112496 181432 112502 181484
rect 112438 180820 112444 180872
rect 112496 180860 112502 180872
rect 163590 180860 163596 180872
rect 112496 180832 163596 180860
rect 112496 180820 112502 180832
rect 163590 180820 163596 180832
rect 163648 180820 163654 180872
rect 71038 180072 71044 180124
rect 71096 180112 71102 180124
rect 167454 180112 167460 180124
rect 71096 180084 167460 180112
rect 71096 180072 71102 180084
rect 167454 180072 167460 180084
rect 167512 180072 167518 180124
rect 97258 177352 97264 177404
rect 97316 177392 97322 177404
rect 123202 177392 123208 177404
rect 97316 177364 123208 177392
rect 97316 177352 97322 177364
rect 123202 177352 123208 177364
rect 123260 177352 123266 177404
rect 68922 177284 68928 177336
rect 68980 177324 68986 177336
rect 167454 177324 167460 177336
rect 68980 177296 167460 177324
rect 68980 177284 68986 177296
rect 167454 177284 167460 177296
rect 167512 177284 167518 177336
rect 123202 176672 123208 176724
rect 123260 176712 123266 176724
rect 123662 176712 123668 176724
rect 123260 176684 123668 176712
rect 123260 176672 123266 176684
rect 123662 176672 123668 176684
rect 123720 176712 123726 176724
rect 166626 176712 166632 176724
rect 123720 176684 166632 176712
rect 123720 176672 123726 176684
rect 166626 176672 166632 176684
rect 166684 176672 166690 176724
rect 65702 175924 65708 175976
rect 65760 175964 65766 175976
rect 69382 175964 69388 175976
rect 65760 175936 69388 175964
rect 65760 175924 65766 175936
rect 69382 175924 69388 175936
rect 69440 175964 69446 175976
rect 168098 175964 168104 175976
rect 69440 175936 168104 175964
rect 69440 175924 69446 175936
rect 168098 175924 168104 175936
rect 168156 175924 168162 175976
rect 233050 175176 233056 175228
rect 233108 175216 233114 175228
rect 494054 175216 494060 175228
rect 233108 175188 494060 175216
rect 233108 175176 233114 175188
rect 494054 175176 494060 175188
rect 494112 175176 494118 175228
rect 111242 174496 111248 174548
rect 111300 174536 111306 174548
rect 140774 174536 140780 174548
rect 111300 174508 140780 174536
rect 111300 174496 111306 174508
rect 140774 174496 140780 174508
rect 140832 174496 140838 174548
rect 140774 173884 140780 173936
rect 140832 173924 140838 173936
rect 141510 173924 141516 173936
rect 140832 173896 141516 173924
rect 140832 173884 140838 173896
rect 141510 173884 141516 173896
rect 141568 173924 141574 173936
rect 168926 173924 168932 173936
rect 141568 173896 168932 173924
rect 141568 173884 141574 173896
rect 168926 173884 168932 173896
rect 168984 173884 168990 173936
rect 80974 173204 80980 173256
rect 81032 173244 81038 173256
rect 114462 173244 114468 173256
rect 81032 173216 114468 173244
rect 81032 173204 81038 173216
rect 114462 173204 114468 173216
rect 114520 173204 114526 173256
rect 66714 173136 66720 173188
rect 66772 173176 66778 173188
rect 168742 173176 168748 173188
rect 66772 173148 168748 173176
rect 66772 173136 66778 173148
rect 168742 173136 168748 173148
rect 168800 173136 168806 173188
rect 170306 173000 170312 173052
rect 170364 173000 170370 173052
rect 170324 172848 170352 173000
rect 170306 172796 170312 172848
rect 170364 172796 170370 172848
rect 113910 172524 113916 172576
rect 113968 172564 113974 172576
rect 114462 172564 114468 172576
rect 113968 172536 114468 172564
rect 113968 172524 113974 172536
rect 114462 172524 114468 172536
rect 114520 172564 114526 172576
rect 168742 172564 168748 172576
rect 114520 172536 168748 172564
rect 114520 172524 114526 172536
rect 168742 172524 168748 172536
rect 168800 172524 168806 172576
rect 68646 172456 68652 172508
rect 68704 172496 68710 172508
rect 168098 172496 168104 172508
rect 68704 172468 168104 172496
rect 68704 172456 68710 172468
rect 168098 172456 168104 172468
rect 168156 172456 168162 172508
rect 112530 171912 112536 171964
rect 112588 171952 112594 171964
rect 123754 171952 123760 171964
rect 112588 171924 123760 171952
rect 112588 171912 112594 171924
rect 123754 171912 123760 171924
rect 123812 171912 123818 171964
rect 111150 171844 111156 171896
rect 111208 171884 111214 171896
rect 134702 171884 134708 171896
rect 111208 171856 134708 171884
rect 111208 171844 111214 171856
rect 134702 171844 134708 171856
rect 134760 171844 134766 171896
rect 70486 171776 70492 171828
rect 70544 171816 70550 171828
rect 170398 171816 170404 171828
rect 70544 171788 170404 171816
rect 70544 171776 70550 171788
rect 170398 171776 170404 171788
rect 170456 171776 170462 171828
rect 231762 171776 231768 171828
rect 231820 171816 231826 171828
rect 462314 171816 462320 171828
rect 231820 171788 462320 171816
rect 231820 171776 231826 171788
rect 462314 171776 462320 171788
rect 462372 171776 462378 171828
rect 134702 171164 134708 171216
rect 134760 171204 134766 171216
rect 169846 171204 169852 171216
rect 134760 171176 169852 171204
rect 134760 171164 134766 171176
rect 169846 171164 169852 171176
rect 169904 171164 169910 171216
rect 123754 171096 123760 171148
rect 123812 171136 123818 171148
rect 169570 171136 169576 171148
rect 123812 171108 169576 171136
rect 123812 171096 123818 171108
rect 169570 171096 169576 171108
rect 169628 171096 169634 171148
rect 231670 171028 231676 171080
rect 231728 171068 231734 171080
rect 231946 171068 231952 171080
rect 231728 171040 231952 171068
rect 231728 171028 231734 171040
rect 231946 171028 231952 171040
rect 232004 171028 232010 171080
rect 170490 170824 170496 170876
rect 170548 170824 170554 170876
rect 170508 170672 170536 170824
rect 96430 170620 96436 170672
rect 96488 170660 96494 170672
rect 125594 170660 125600 170672
rect 96488 170632 125600 170660
rect 96488 170620 96494 170632
rect 125594 170620 125600 170632
rect 125652 170660 125658 170672
rect 126882 170660 126888 170672
rect 125652 170632 126888 170660
rect 125652 170620 125658 170632
rect 126882 170620 126888 170632
rect 126940 170620 126946 170672
rect 170490 170620 170496 170672
rect 170548 170620 170554 170672
rect 83550 170552 83556 170604
rect 83608 170592 83614 170604
rect 115382 170592 115388 170604
rect 83608 170564 115388 170592
rect 83608 170552 83614 170564
rect 115382 170552 115388 170564
rect 115440 170552 115446 170604
rect 169846 170552 169852 170604
rect 169904 170552 169910 170604
rect 109310 170484 109316 170536
rect 109368 170524 109374 170536
rect 143442 170524 143448 170536
rect 109368 170496 143448 170524
rect 109368 170484 109374 170496
rect 143442 170484 143448 170496
rect 143500 170484 143506 170536
rect 75178 170416 75184 170468
rect 75236 170456 75242 170468
rect 109218 170456 109224 170468
rect 75236 170428 109224 170456
rect 75236 170416 75242 170428
rect 109218 170416 109224 170428
rect 109276 170416 109282 170468
rect 169864 170400 169892 170552
rect 69290 170348 69296 170400
rect 69348 170388 69354 170400
rect 168098 170388 168104 170400
rect 69348 170360 168104 170388
rect 69348 170348 69354 170360
rect 168098 170348 168104 170360
rect 168156 170348 168162 170400
rect 169846 170348 169852 170400
rect 169904 170348 169910 170400
rect 228818 170348 228824 170400
rect 228876 170388 228882 170400
rect 231854 170388 231860 170400
rect 228876 170360 231860 170388
rect 228876 170348 228882 170360
rect 231854 170348 231860 170360
rect 231912 170348 231918 170400
rect 168650 170280 168656 170332
rect 168708 170320 168714 170332
rect 173250 170320 173256 170332
rect 168708 170292 173256 170320
rect 168708 170280 168714 170292
rect 173250 170280 173256 170292
rect 173308 170280 173314 170332
rect 167914 170212 167920 170264
rect 167972 170252 167978 170264
rect 171962 170252 171968 170264
rect 167972 170224 171968 170252
rect 167972 170212 167978 170224
rect 171962 170212 171968 170224
rect 172020 170212 172026 170264
rect 173894 170212 173900 170264
rect 173952 170212 173958 170264
rect 175182 170212 175188 170264
rect 175240 170212 175246 170264
rect 176470 170252 176476 170264
rect 175292 170224 176476 170252
rect 170398 170184 170404 170196
rect 161446 170156 170404 170184
rect 142982 169940 142988 169992
rect 143040 169980 143046 169992
rect 143442 169980 143448 169992
rect 143040 169952 143448 169980
rect 143040 169940 143046 169952
rect 143442 169940 143448 169952
rect 143500 169980 143506 169992
rect 161446 169980 161474 170156
rect 170398 170144 170404 170156
rect 170456 170144 170462 170196
rect 170030 170048 170036 170060
rect 143500 169952 161474 169980
rect 166000 170020 170036 170048
rect 143500 169940 143506 169952
rect 126882 169872 126888 169924
rect 126940 169912 126946 169924
rect 166000 169912 166028 170020
rect 170030 170008 170036 170020
rect 170088 170008 170094 170060
rect 173912 169992 173940 170212
rect 175200 169992 175228 170212
rect 175292 169992 175320 170224
rect 176470 170212 176476 170224
rect 176528 170212 176534 170264
rect 177758 170212 177764 170264
rect 177816 170212 177822 170264
rect 178402 170212 178408 170264
rect 178460 170212 178466 170264
rect 179690 170212 179696 170264
rect 179748 170212 179754 170264
rect 180978 170212 180984 170264
rect 181036 170212 181042 170264
rect 181622 170212 181628 170264
rect 181680 170212 181686 170264
rect 182910 170212 182916 170264
rect 182968 170212 182974 170264
rect 184198 170212 184204 170264
rect 184256 170212 184262 170264
rect 185486 170212 185492 170264
rect 185544 170212 185550 170264
rect 186130 170212 186136 170264
rect 186188 170212 186194 170264
rect 187418 170212 187424 170264
rect 187476 170212 187482 170264
rect 188706 170212 188712 170264
rect 188764 170212 188770 170264
rect 189350 170212 189356 170264
rect 189408 170212 189414 170264
rect 190638 170252 190644 170264
rect 189460 170224 190644 170252
rect 177776 169992 177804 170212
rect 178420 169992 178448 170212
rect 179708 169992 179736 170212
rect 180996 169992 181024 170212
rect 181640 169992 181668 170212
rect 182928 169992 182956 170212
rect 184216 169992 184244 170212
rect 185504 169992 185532 170212
rect 186148 169992 186176 170212
rect 187436 169992 187464 170212
rect 188724 169992 188752 170212
rect 189368 169992 189396 170212
rect 189460 169992 189488 170224
rect 190638 170212 190644 170224
rect 190696 170212 190702 170264
rect 191926 170212 191932 170264
rect 191984 170212 191990 170264
rect 193214 170212 193220 170264
rect 193272 170212 193278 170264
rect 193858 170212 193864 170264
rect 193916 170212 193922 170264
rect 195146 170212 195152 170264
rect 195204 170212 195210 170264
rect 196434 170212 196440 170264
rect 196492 170212 196498 170264
rect 197078 170252 197084 170264
rect 196544 170224 197084 170252
rect 191944 169992 191972 170212
rect 193232 169992 193260 170212
rect 193876 169992 193904 170212
rect 195164 169992 195192 170212
rect 196452 169992 196480 170212
rect 196544 169992 196572 170224
rect 197078 170212 197084 170224
rect 197136 170212 197142 170264
rect 198366 170212 198372 170264
rect 198424 170212 198430 170264
rect 199654 170212 199660 170264
rect 199712 170212 199718 170264
rect 200942 170212 200948 170264
rect 201000 170252 201006 170264
rect 201000 170224 201448 170252
rect 201000 170212 201006 170224
rect 198384 169992 198412 170212
rect 199672 169992 199700 170212
rect 201420 169992 201448 170224
rect 201586 170212 201592 170264
rect 201644 170212 201650 170264
rect 202874 170212 202880 170264
rect 202932 170212 202938 170264
rect 204162 170212 204168 170264
rect 204220 170212 204226 170264
rect 204806 170212 204812 170264
rect 204864 170212 204870 170264
rect 206094 170212 206100 170264
rect 206152 170212 206158 170264
rect 207382 170212 207388 170264
rect 207440 170212 207446 170264
rect 208670 170212 208676 170264
rect 208728 170212 208734 170264
rect 209314 170212 209320 170264
rect 209372 170212 209378 170264
rect 210602 170212 210608 170264
rect 210660 170212 210666 170264
rect 211890 170212 211896 170264
rect 211948 170212 211954 170264
rect 212534 170212 212540 170264
rect 212592 170212 212598 170264
rect 213822 170212 213828 170264
rect 213880 170212 213886 170264
rect 215110 170212 215116 170264
rect 215168 170212 215174 170264
rect 216398 170212 216404 170264
rect 216456 170212 216462 170264
rect 217042 170212 217048 170264
rect 217100 170212 217106 170264
rect 218330 170212 218336 170264
rect 218388 170212 218394 170264
rect 219618 170212 219624 170264
rect 219676 170212 219682 170264
rect 220262 170212 220268 170264
rect 220320 170212 220326 170264
rect 221550 170212 221556 170264
rect 221608 170212 221614 170264
rect 222838 170212 222844 170264
rect 222896 170212 222902 170264
rect 224126 170212 224132 170264
rect 224184 170212 224190 170264
rect 224770 170212 224776 170264
rect 224828 170212 224834 170264
rect 226058 170212 226064 170264
rect 226116 170212 226122 170264
rect 227346 170212 227352 170264
rect 227404 170212 227410 170264
rect 201604 169992 201632 170212
rect 202892 169992 202920 170212
rect 204180 169992 204208 170212
rect 204824 169992 204852 170212
rect 206112 169992 206140 170212
rect 207400 169992 207428 170212
rect 208688 169992 208716 170212
rect 173894 169940 173900 169992
rect 173952 169940 173958 169992
rect 175182 169940 175188 169992
rect 175240 169940 175246 169992
rect 175274 169940 175280 169992
rect 175332 169940 175338 169992
rect 177758 169940 177764 169992
rect 177816 169940 177822 169992
rect 178402 169940 178408 169992
rect 178460 169940 178466 169992
rect 179690 169940 179696 169992
rect 179748 169940 179754 169992
rect 180978 169940 180984 169992
rect 181036 169940 181042 169992
rect 181622 169940 181628 169992
rect 181680 169940 181686 169992
rect 182910 169940 182916 169992
rect 182968 169940 182974 169992
rect 184198 169940 184204 169992
rect 184256 169940 184262 169992
rect 185486 169940 185492 169992
rect 185544 169940 185550 169992
rect 186130 169940 186136 169992
rect 186188 169940 186194 169992
rect 187418 169940 187424 169992
rect 187476 169940 187482 169992
rect 188706 169940 188712 169992
rect 188764 169940 188770 169992
rect 189350 169940 189356 169992
rect 189408 169940 189414 169992
rect 189442 169940 189448 169992
rect 189500 169940 189506 169992
rect 191926 169940 191932 169992
rect 191984 169940 191990 169992
rect 193214 169940 193220 169992
rect 193272 169940 193278 169992
rect 193858 169940 193864 169992
rect 193916 169940 193922 169992
rect 195146 169940 195152 169992
rect 195204 169940 195210 169992
rect 196434 169940 196440 169992
rect 196492 169940 196498 169992
rect 196526 169940 196532 169992
rect 196584 169940 196590 169992
rect 198366 169940 198372 169992
rect 198424 169940 198430 169992
rect 199654 169940 199660 169992
rect 199712 169940 199718 169992
rect 201402 169940 201408 169992
rect 201460 169940 201466 169992
rect 201586 169940 201592 169992
rect 201644 169940 201650 169992
rect 202874 169940 202880 169992
rect 202932 169940 202938 169992
rect 204162 169940 204168 169992
rect 204220 169940 204226 169992
rect 204806 169940 204812 169992
rect 204864 169940 204870 169992
rect 206094 169940 206100 169992
rect 206152 169940 206158 169992
rect 207382 169940 207388 169992
rect 207440 169940 207446 169992
rect 208670 169940 208676 169992
rect 208728 169940 208734 169992
rect 170950 169912 170956 169924
rect 126940 169884 166028 169912
rect 166184 169884 170956 169912
rect 126940 169872 126946 169884
rect 115382 169804 115388 169856
rect 115440 169844 115446 169856
rect 166184 169844 166212 169884
rect 170950 169872 170956 169884
rect 171008 169872 171014 169924
rect 171042 169844 171048 169856
rect 115440 169816 166212 169844
rect 166276 169816 171048 169844
rect 115440 169804 115446 169816
rect 109218 169736 109224 169788
rect 109276 169776 109282 169788
rect 109678 169776 109684 169788
rect 109276 169748 109684 169776
rect 109276 169736 109282 169748
rect 109678 169736 109684 169748
rect 109736 169776 109742 169788
rect 166276 169776 166304 169816
rect 171042 169804 171048 169816
rect 171100 169804 171106 169856
rect 109736 169748 166304 169776
rect 109736 169736 109742 169748
rect 168006 169736 168012 169788
rect 168064 169776 168070 169788
rect 169662 169776 169668 169788
rect 168064 169748 169668 169776
rect 168064 169736 168070 169748
rect 169662 169736 169668 169748
rect 169720 169736 169726 169788
rect 166442 169668 166448 169720
rect 166500 169708 166506 169720
rect 209332 169708 209360 170212
rect 210620 169992 210648 170212
rect 211908 169992 211936 170212
rect 212552 169992 212580 170212
rect 213840 169992 213868 170212
rect 215128 169992 215156 170212
rect 216416 169992 216444 170212
rect 217060 169992 217088 170212
rect 218348 169992 218376 170212
rect 219636 169992 219664 170212
rect 220280 169992 220308 170212
rect 221568 169992 221596 170212
rect 222856 169992 222884 170212
rect 210602 169940 210608 169992
rect 210660 169940 210666 169992
rect 211890 169940 211896 169992
rect 211948 169940 211954 169992
rect 212534 169940 212540 169992
rect 212592 169940 212598 169992
rect 213822 169940 213828 169992
rect 213880 169940 213886 169992
rect 215110 169940 215116 169992
rect 215168 169940 215174 169992
rect 216398 169940 216404 169992
rect 216456 169940 216462 169992
rect 217042 169940 217048 169992
rect 217100 169940 217106 169992
rect 218330 169940 218336 169992
rect 218388 169940 218394 169992
rect 219618 169940 219624 169992
rect 219676 169940 219682 169992
rect 220262 169940 220268 169992
rect 220320 169940 220326 169992
rect 221550 169940 221556 169992
rect 221608 169940 221614 169992
rect 222838 169940 222844 169992
rect 222896 169940 222902 169992
rect 224144 169708 224172 170212
rect 224788 169992 224816 170212
rect 226076 169992 226104 170212
rect 227364 169992 227392 170212
rect 224770 169940 224776 169992
rect 224828 169940 224834 169992
rect 226058 169940 226064 169992
rect 226116 169940 226122 169992
rect 227346 169940 227352 169992
rect 227404 169940 227410 169992
rect 166500 169680 209360 169708
rect 215266 169680 224172 169708
rect 166500 169668 166506 169680
rect 115290 169600 115296 169652
rect 115348 169640 115354 169652
rect 215266 169640 215294 169680
rect 115348 169612 215294 169640
rect 115348 169600 115354 169612
rect 108298 169572 108304 169584
rect 103486 169544 108304 169572
rect 73246 169328 73252 169380
rect 73304 169368 73310 169380
rect 103486 169368 103514 169544
rect 108298 169532 108304 169544
rect 108356 169572 108362 169584
rect 173894 169572 173900 169584
rect 108356 169544 173900 169572
rect 108356 169532 108362 169544
rect 173894 169532 173900 169544
rect 173952 169532 173958 169584
rect 175182 169532 175188 169584
rect 175240 169572 175246 169584
rect 238018 169572 238024 169584
rect 175240 169544 238024 169572
rect 175240 169532 175246 169544
rect 238018 169532 238024 169544
rect 238076 169532 238082 169584
rect 166350 169464 166356 169516
rect 166408 169504 166414 169516
rect 215110 169504 215116 169516
rect 166408 169476 215116 169504
rect 166408 169464 166414 169476
rect 215110 169464 215116 169476
rect 215168 169464 215174 169516
rect 118050 169396 118056 169448
rect 118108 169436 118114 169448
rect 181162 169436 181168 169448
rect 118108 169408 181168 169436
rect 118108 169396 118114 169408
rect 181162 169396 181168 169408
rect 181220 169396 181226 169448
rect 198366 169396 198372 169448
rect 198424 169436 198430 169448
rect 235258 169436 235264 169448
rect 198424 169408 235264 169436
rect 198424 169396 198430 169408
rect 235258 169396 235264 169408
rect 235316 169396 235322 169448
rect 73304 169340 103514 169368
rect 73304 169328 73310 169340
rect 170490 169328 170496 169380
rect 170548 169368 170554 169380
rect 213822 169368 213828 169380
rect 170548 169340 213828 169368
rect 170548 169328 170554 169340
rect 213822 169328 213828 169340
rect 213880 169328 213886 169380
rect 79318 169260 79324 169312
rect 79376 169300 79382 169312
rect 110690 169300 110696 169312
rect 79376 169272 110696 169300
rect 79376 169260 79382 169272
rect 110690 169260 110696 169272
rect 110748 169260 110754 169312
rect 170214 169260 170220 169312
rect 170272 169300 170278 169312
rect 207382 169300 207388 169312
rect 170272 169272 207388 169300
rect 170272 169260 170278 169272
rect 207382 169260 207388 169272
rect 207440 169260 207446 169312
rect 94590 169192 94596 169244
rect 94648 169232 94654 169244
rect 127802 169232 127808 169244
rect 94648 169204 127808 169232
rect 94648 169192 94654 169204
rect 127802 169192 127808 169204
rect 127860 169232 127866 169244
rect 196526 169232 196532 169244
rect 127860 169204 196532 169232
rect 127860 169192 127866 169204
rect 196526 169192 196532 169204
rect 196584 169192 196590 169244
rect 87598 169124 87604 169176
rect 87656 169164 87662 169176
rect 122098 169164 122104 169176
rect 87656 169136 122104 169164
rect 87656 169124 87662 169136
rect 122098 169124 122104 169136
rect 122156 169164 122162 169176
rect 189442 169164 189448 169176
rect 122156 169136 189448 169164
rect 122156 169124 122162 169136
rect 189442 169124 189448 169136
rect 189500 169124 189506 169176
rect 84194 169056 84200 169108
rect 84252 169096 84258 169108
rect 156690 169096 156696 169108
rect 84252 169068 156696 169096
rect 84252 169056 84258 169068
rect 156690 169056 156696 169068
rect 156748 169056 156754 169108
rect 169018 169056 169024 169108
rect 169076 169096 169082 169108
rect 229278 169096 229284 169108
rect 169076 169068 229284 169096
rect 169076 169056 169082 169068
rect 229278 169056 229284 169068
rect 229336 169056 229342 169108
rect 103422 168988 103428 169040
rect 103480 169028 103486 169040
rect 133322 169028 133328 169040
rect 103480 169000 133328 169028
rect 103480 168988 103486 169000
rect 133322 168988 133328 169000
rect 133380 169028 133386 169040
rect 208670 169028 208676 169040
rect 133380 169000 208676 169028
rect 133380 168988 133386 169000
rect 208670 168988 208676 169000
rect 208728 168988 208734 169040
rect 209682 168988 209688 169040
rect 209740 169028 209746 169040
rect 580442 169028 580448 169040
rect 209740 169000 580448 169028
rect 209740 168988 209746 169000
rect 580442 168988 580448 169000
rect 580500 168988 580506 169040
rect 166258 168920 166264 168972
rect 166316 168960 166322 168972
rect 201402 168960 201408 168972
rect 166316 168932 201408 168960
rect 166316 168920 166322 168932
rect 201402 168920 201408 168932
rect 201460 168920 201466 168972
rect 110690 168852 110696 168904
rect 110748 168892 110754 168904
rect 111150 168892 111156 168904
rect 110748 168864 111156 168892
rect 110748 168852 110754 168864
rect 111150 168852 111156 168864
rect 111208 168892 111214 168904
rect 178402 168892 178408 168904
rect 111208 168864 178408 168892
rect 111208 168852 111214 168864
rect 178402 168852 178408 168864
rect 178460 168852 178466 168904
rect 184934 168852 184940 168904
rect 184992 168892 184998 168904
rect 186130 168892 186136 168904
rect 184992 168864 186136 168892
rect 184992 168852 184998 168864
rect 186130 168852 186136 168864
rect 186188 168892 186194 168904
rect 396718 168892 396724 168904
rect 186188 168864 396724 168892
rect 186188 168852 186194 168864
rect 396718 168852 396724 168864
rect 396776 168852 396782 168904
rect 156690 168376 156696 168428
rect 156748 168416 156754 168428
rect 187418 168416 187424 168428
rect 156748 168388 187424 168416
rect 156748 168376 156754 168388
rect 187418 168376 187424 168388
rect 187476 168376 187482 168428
rect 171042 168308 171048 168360
rect 171100 168348 171106 168360
rect 175274 168348 175280 168360
rect 171100 168320 175280 168348
rect 171100 168308 171106 168320
rect 175274 168308 175280 168320
rect 175332 168308 175338 168360
rect 196434 168308 196440 168360
rect 196492 168348 196498 168360
rect 203426 168348 203432 168360
rect 196492 168320 203432 168348
rect 196492 168308 196498 168320
rect 203426 168308 203432 168320
rect 203484 168308 203490 168360
rect 226058 168308 226064 168360
rect 226116 168348 226122 168360
rect 347774 168348 347780 168360
rect 226116 168320 347780 168348
rect 226116 168308 226122 168320
rect 347774 168308 347780 168320
rect 347832 168308 347838 168360
rect 123846 168240 123852 168292
rect 123904 168280 123910 168292
rect 228726 168280 228732 168292
rect 123904 168252 228732 168280
rect 123904 168240 123910 168252
rect 228726 168240 228732 168252
rect 228784 168240 228790 168292
rect 169570 168172 169576 168224
rect 169628 168212 169634 168224
rect 220262 168212 220268 168224
rect 169628 168184 220268 168212
rect 169628 168172 169634 168184
rect 220262 168172 220268 168184
rect 220320 168172 220326 168224
rect 221550 168172 221556 168224
rect 221608 168212 221614 168224
rect 299474 168212 299480 168224
rect 221608 168184 299480 168212
rect 221608 168172 221614 168184
rect 299474 168172 299480 168184
rect 299532 168172 299538 168224
rect 166626 168104 166632 168156
rect 166684 168144 166690 168156
rect 202874 168144 202880 168156
rect 166684 168116 202880 168144
rect 166684 168104 166690 168116
rect 202874 168104 202880 168116
rect 202932 168104 202938 168156
rect 218330 168104 218336 168156
rect 218388 168144 218394 168156
rect 239398 168144 239404 168156
rect 218388 168116 239404 168144
rect 218388 168104 218394 168116
rect 239398 168104 239404 168116
rect 239456 168104 239462 168156
rect 169846 168036 169852 168088
rect 169904 168076 169910 168088
rect 219618 168076 219624 168088
rect 169904 168048 219624 168076
rect 169904 168036 169910 168048
rect 219618 168036 219624 168048
rect 219676 168036 219682 168088
rect 170398 167968 170404 168020
rect 170456 168008 170462 168020
rect 217042 168008 217048 168020
rect 170456 167980 217048 168008
rect 170456 167968 170462 167980
rect 217042 167968 217048 167980
rect 217100 167968 217106 168020
rect 181162 167900 181168 167952
rect 181220 167940 181226 167952
rect 227346 167940 227352 167952
rect 181220 167912 227352 167940
rect 181220 167900 181226 167912
rect 227346 167900 227352 167912
rect 227404 167900 227410 167952
rect 170030 167832 170036 167884
rect 170088 167872 170094 167884
rect 201586 167872 201592 167884
rect 170088 167844 201592 167872
rect 170088 167832 170094 167844
rect 201586 167832 201592 167844
rect 201644 167832 201650 167884
rect 163498 167764 163504 167816
rect 163556 167804 163562 167816
rect 195146 167804 195152 167816
rect 163556 167776 195152 167804
rect 163556 167764 163562 167776
rect 195146 167764 195152 167776
rect 195204 167764 195210 167816
rect 163958 167696 163964 167748
rect 164016 167736 164022 167748
rect 168650 167736 168656 167748
rect 164016 167708 168656 167736
rect 164016 167696 164022 167708
rect 168650 167696 168656 167708
rect 168708 167696 168714 167748
rect 195238 167696 195244 167748
rect 195296 167736 195302 167748
rect 233234 167736 233240 167748
rect 195296 167708 233240 167736
rect 195296 167696 195302 167708
rect 233234 167696 233240 167708
rect 233292 167696 233298 167748
rect 86218 167628 86224 167680
rect 86276 167668 86282 167680
rect 111242 167668 111248 167680
rect 86276 167640 111248 167668
rect 86276 167628 86282 167640
rect 111242 167628 111248 167640
rect 111300 167668 111306 167680
rect 177758 167668 177764 167680
rect 111300 167640 177764 167668
rect 111300 167628 111306 167640
rect 177758 167628 177764 167640
rect 177816 167628 177822 167680
rect 195330 167628 195336 167680
rect 195388 167668 195394 167680
rect 234706 167668 234712 167680
rect 195388 167640 234712 167668
rect 195388 167628 195394 167640
rect 234706 167628 234712 167640
rect 234764 167628 234770 167680
rect 164050 167560 164056 167612
rect 164108 167600 164114 167612
rect 167914 167600 167920 167612
rect 164108 167572 167920 167600
rect 164108 167560 164114 167572
rect 167914 167560 167920 167572
rect 167972 167560 167978 167612
rect 189350 167560 189356 167612
rect 189408 167600 189414 167612
rect 204346 167600 204352 167612
rect 189408 167572 204352 167600
rect 189408 167560 189414 167572
rect 204346 167560 204352 167572
rect 204404 167560 204410 167612
rect 162394 167492 162400 167544
rect 162452 167532 162458 167544
rect 224770 167532 224776 167544
rect 162452 167504 224776 167532
rect 162452 167492 162458 167504
rect 224770 167492 224776 167504
rect 224828 167492 224834 167544
rect 163590 167424 163596 167476
rect 163648 167464 163654 167476
rect 179690 167464 179696 167476
rect 163648 167436 179696 167464
rect 163648 167424 163654 167436
rect 179690 167424 179696 167436
rect 179748 167424 179754 167476
rect 193214 167424 193220 167476
rect 193272 167464 193278 167476
rect 244918 167464 244924 167476
rect 193272 167436 244924 167464
rect 193272 167424 193278 167436
rect 244918 167424 244924 167436
rect 244976 167424 244982 167476
rect 156874 167356 156880 167408
rect 156932 167396 156938 167408
rect 185486 167396 185492 167408
rect 156932 167368 185492 167396
rect 156932 167356 156938 167368
rect 185486 167356 185492 167368
rect 185544 167356 185550 167408
rect 182910 167288 182916 167340
rect 182968 167328 182974 167340
rect 209682 167328 209688 167340
rect 182968 167300 209688 167328
rect 182968 167288 182974 167300
rect 209682 167288 209688 167300
rect 209740 167288 209746 167340
rect 548518 166948 548524 167000
rect 548576 166988 548582 167000
rect 580166 166988 580172 167000
rect 548576 166960 580172 166988
rect 548576 166948 548582 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 226978 166404 226984 166456
rect 227036 166444 227042 166456
rect 232222 166444 232228 166456
rect 227036 166416 232228 166444
rect 227036 166404 227042 166416
rect 232222 166404 232228 166416
rect 232280 166404 232286 166456
rect 215202 166336 215208 166388
rect 215260 166376 215266 166388
rect 232498 166376 232504 166388
rect 215260 166348 232504 166376
rect 215260 166336 215266 166348
rect 232498 166336 232504 166348
rect 232556 166336 232562 166388
rect 202230 166268 202236 166320
rect 202288 166308 202294 166320
rect 230014 166308 230020 166320
rect 202288 166280 230020 166308
rect 202288 166268 202294 166280
rect 230014 166268 230020 166280
rect 230072 166268 230078 166320
rect 108482 165520 108488 165572
rect 108540 165560 108546 165572
rect 233418 165560 233424 165572
rect 108540 165532 233424 165560
rect 108540 165520 108546 165532
rect 233418 165520 233424 165532
rect 233476 165520 233482 165572
rect 108850 165452 108856 165504
rect 108908 165492 108914 165504
rect 232406 165492 232412 165504
rect 108908 165464 232412 165492
rect 108908 165452 108914 165464
rect 232406 165452 232412 165464
rect 232464 165452 232470 165504
rect 108758 165384 108764 165436
rect 108816 165424 108822 165436
rect 229554 165424 229560 165436
rect 108816 165396 229560 165424
rect 108816 165384 108822 165396
rect 229554 165384 229560 165396
rect 229612 165384 229618 165436
rect 120994 165316 121000 165368
rect 121052 165356 121058 165368
rect 229370 165356 229376 165368
rect 121052 165328 229376 165356
rect 121052 165316 121058 165328
rect 229370 165316 229376 165328
rect 229428 165316 229434 165368
rect 124398 165288 124404 165300
rect 122806 165260 124404 165288
rect 111702 164908 111708 164960
rect 111760 164948 111766 164960
rect 122806 164948 122834 165260
rect 124398 165248 124404 165260
rect 124456 165288 124462 165300
rect 231854 165288 231860 165300
rect 124456 165260 231860 165288
rect 124456 165248 124462 165260
rect 231854 165248 231860 165260
rect 231912 165248 231918 165300
rect 144270 165180 144276 165232
rect 144328 165220 144334 165232
rect 144822 165220 144828 165232
rect 144328 165192 144828 165220
rect 144328 165180 144334 165192
rect 144822 165180 144828 165192
rect 144880 165220 144886 165232
rect 233510 165220 233516 165232
rect 144880 165192 233516 165220
rect 144880 165180 144886 165192
rect 233510 165180 233516 165192
rect 233568 165180 233574 165232
rect 148410 165112 148416 165164
rect 148468 165152 148474 165164
rect 148962 165152 148968 165164
rect 148468 165124 148968 165152
rect 148468 165112 148474 165124
rect 148962 165112 148968 165124
rect 149020 165152 149026 165164
rect 232774 165152 232780 165164
rect 149020 165124 232780 165152
rect 149020 165112 149026 165124
rect 232774 165112 232780 165124
rect 232832 165112 232838 165164
rect 152550 165044 152556 165096
rect 152608 165084 152614 165096
rect 153102 165084 153108 165096
rect 152608 165056 153108 165084
rect 152608 165044 152614 165056
rect 153102 165044 153108 165056
rect 153160 165084 153166 165096
rect 231946 165084 231952 165096
rect 153160 165056 231952 165084
rect 153160 165044 153166 165056
rect 231946 165044 231952 165056
rect 232004 165044 232010 165096
rect 164878 164976 164884 165028
rect 164936 165016 164942 165028
rect 188706 165016 188712 165028
rect 164936 164988 188712 165016
rect 164936 164976 164942 164988
rect 188706 164976 188712 164988
rect 188764 164976 188770 165028
rect 209038 164976 209044 165028
rect 209096 165016 209102 165028
rect 232682 165016 232688 165028
rect 209096 164988 232688 165016
rect 209096 164976 209102 164988
rect 232682 164976 232688 164988
rect 232740 164976 232746 165028
rect 111760 164920 122834 164948
rect 111760 164908 111766 164920
rect 166350 164908 166356 164960
rect 166408 164948 166414 164960
rect 193858 164948 193864 164960
rect 166408 164920 193864 164948
rect 166408 164908 166414 164920
rect 193858 164908 193864 164920
rect 193916 164908 193922 164960
rect 202138 164908 202144 164960
rect 202196 164948 202202 164960
rect 230934 164948 230940 164960
rect 202196 164920 230940 164948
rect 202196 164908 202202 164920
rect 230934 164908 230940 164920
rect 230992 164908 230998 164960
rect 119338 164840 119344 164892
rect 119396 164880 119402 164892
rect 229462 164880 229468 164892
rect 119396 164852 229468 164880
rect 119396 164840 119402 164852
rect 229462 164840 229468 164852
rect 229520 164840 229526 164892
rect 166258 164772 166264 164824
rect 166316 164812 166322 164824
rect 184198 164812 184204 164824
rect 166316 164784 184204 164812
rect 166316 164772 166322 164784
rect 184198 164772 184204 164784
rect 184256 164772 184262 164824
rect 163774 164704 163780 164756
rect 163832 164744 163838 164756
rect 180978 164744 180984 164756
rect 163832 164716 180984 164744
rect 163832 164704 163838 164716
rect 180978 164704 180984 164716
rect 181036 164704 181042 164756
rect 163866 164636 163872 164688
rect 163924 164676 163930 164688
rect 181622 164676 181628 164688
rect 163924 164648 181628 164676
rect 163924 164636 163930 164648
rect 181622 164636 181628 164648
rect 181680 164636 181686 164688
rect 224862 163548 224868 163600
rect 224920 163588 224926 163600
rect 232038 163588 232044 163600
rect 224920 163560 232044 163588
rect 224920 163548 224926 163560
rect 232038 163548 232044 163560
rect 232096 163548 232102 163600
rect 164970 163480 164976 163532
rect 165028 163520 165034 163532
rect 201494 163520 201500 163532
rect 165028 163492 201500 163520
rect 165028 163480 165034 163492
rect 201494 163480 201500 163492
rect 201552 163520 201558 163532
rect 231026 163520 231032 163532
rect 201552 163492 231032 163520
rect 201552 163480 201558 163492
rect 231026 163480 231032 163492
rect 231084 163480 231090 163532
rect 166718 162120 166724 162172
rect 166776 162160 166782 162172
rect 191926 162160 191932 162172
rect 166776 162132 191932 162160
rect 166776 162120 166782 162132
rect 191926 162120 191932 162132
rect 191984 162120 191990 162172
rect 201402 162120 201408 162172
rect 201460 162160 201466 162172
rect 580258 162160 580264 162172
rect 201460 162132 580264 162160
rect 201460 162120 201466 162132
rect 580258 162120 580264 162132
rect 580316 162120 580322 162172
rect 199930 160692 199936 160744
rect 199988 160732 199994 160744
rect 230842 160732 230848 160744
rect 199988 160704 230848 160732
rect 199988 160692 199994 160704
rect 230842 160692 230848 160704
rect 230900 160692 230906 160744
rect 217962 159332 217968 159384
rect 218020 159372 218026 159384
rect 229094 159372 229100 159384
rect 218020 159344 229100 159372
rect 218020 159332 218026 159344
rect 229094 159332 229100 159344
rect 229152 159332 229158 159384
rect 2958 149064 2964 149116
rect 3016 149104 3022 149116
rect 106458 149104 106464 149116
rect 3016 149076 106464 149104
rect 3016 149064 3022 149076
rect 106458 149064 106464 149076
rect 106516 149064 106522 149116
rect 202322 142808 202328 142860
rect 202380 142848 202386 142860
rect 231302 142848 231308 142860
rect 202380 142820 231308 142848
rect 202380 142808 202386 142820
rect 231302 142808 231308 142820
rect 231360 142808 231366 142860
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 61746 137952 61752 137964
rect 3568 137924 61752 137952
rect 3568 137912 3574 137924
rect 61746 137912 61752 137924
rect 61804 137952 61810 137964
rect 65518 137952 65524 137964
rect 61804 137924 65524 137952
rect 61804 137912 61810 137924
rect 65518 137912 65524 137924
rect 65576 137912 65582 137964
rect 220722 131724 220728 131776
rect 220780 131764 220786 131776
rect 232590 131764 232596 131776
rect 220780 131736 232596 131764
rect 220780 131724 220786 131736
rect 232590 131724 232596 131736
rect 232648 131724 232654 131776
rect 201586 130404 201592 130416
rect 122806 130376 201592 130404
rect 119062 130228 119068 130280
rect 119120 130268 119126 130280
rect 119614 130268 119620 130280
rect 119120 130240 119620 130268
rect 119120 130228 119126 130240
rect 119614 130228 119620 130240
rect 119672 130268 119678 130280
rect 122806 130268 122834 130376
rect 201586 130364 201592 130376
rect 201644 130404 201650 130416
rect 202230 130404 202236 130416
rect 201644 130376 202236 130404
rect 201644 130364 201650 130376
rect 202230 130364 202236 130376
rect 202288 130364 202294 130416
rect 119672 130240 122834 130268
rect 119672 130228 119678 130240
rect 122282 129004 122288 129056
rect 122340 129044 122346 129056
rect 219434 129044 219440 129056
rect 122340 129016 219440 129044
rect 122340 129004 122346 129016
rect 219434 129004 219440 129016
rect 219492 129044 219498 129056
rect 220722 129044 220728 129056
rect 219492 129016 220728 129044
rect 219492 129004 219498 129016
rect 220722 129004 220728 129016
rect 220780 129004 220786 129056
rect 169662 127576 169668 127628
rect 169720 127616 169726 127628
rect 580258 127616 580264 127628
rect 169720 127588 580264 127616
rect 169720 127576 169726 127588
rect 580258 127576 580264 127588
rect 580316 127576 580322 127628
rect 234614 126896 234620 126948
rect 234672 126936 234678 126948
rect 580166 126936 580172 126948
rect 234672 126908 580172 126936
rect 234672 126896 234678 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 66990 126216 66996 126268
rect 67048 126256 67054 126268
rect 169018 126256 169024 126268
rect 67048 126228 169024 126256
rect 67048 126216 67054 126228
rect 169018 126216 169024 126228
rect 169076 126256 169082 126268
rect 169662 126256 169668 126268
rect 169076 126228 169668 126256
rect 169076 126216 169082 126228
rect 169662 126216 169668 126228
rect 169720 126216 169726 126268
rect 183554 126216 183560 126268
rect 183612 126256 183618 126268
rect 234614 126256 234620 126268
rect 183612 126228 234620 126256
rect 183612 126216 183618 126228
rect 234614 126216 234620 126228
rect 234672 126216 234678 126268
rect 147030 125468 147036 125520
rect 147088 125508 147094 125520
rect 147582 125508 147588 125520
rect 147088 125480 147588 125508
rect 147088 125468 147094 125480
rect 147582 125468 147588 125480
rect 147640 125468 147646 125520
rect 162486 124992 162492 125044
rect 162544 125032 162550 125044
rect 202230 125032 202236 125044
rect 162544 125004 202236 125032
rect 162544 124992 162550 125004
rect 202230 124992 202236 125004
rect 202288 124992 202294 125044
rect 162578 124924 162584 124976
rect 162636 124964 162642 124976
rect 200482 124964 200488 124976
rect 162636 124936 200488 124964
rect 162636 124924 162642 124936
rect 200482 124924 200488 124936
rect 200540 124924 200546 124976
rect 111610 124856 111616 124908
rect 111668 124896 111674 124908
rect 121454 124896 121460 124908
rect 111668 124868 121460 124896
rect 111668 124856 111674 124868
rect 121454 124856 121460 124868
rect 121512 124856 121518 124908
rect 147030 124856 147036 124908
rect 147088 124896 147094 124908
rect 202046 124896 202052 124908
rect 147088 124868 202052 124896
rect 147088 124856 147094 124868
rect 202046 124856 202052 124868
rect 202104 124856 202110 124908
rect 119890 124788 119896 124840
rect 119948 124828 119954 124840
rect 200022 124828 200028 124840
rect 119948 124800 200028 124828
rect 119948 124788 119954 124800
rect 200022 124788 200028 124800
rect 200080 124788 200086 124840
rect 121362 124720 121368 124772
rect 121420 124760 121426 124772
rect 200390 124760 200396 124772
rect 121420 124732 200396 124760
rect 121420 124720 121426 124732
rect 200390 124720 200396 124732
rect 200448 124720 200454 124772
rect 121086 124652 121092 124704
rect 121144 124692 121150 124704
rect 201770 124692 201776 124704
rect 121144 124664 201776 124692
rect 121144 124652 121150 124664
rect 201770 124652 201776 124664
rect 201828 124652 201834 124704
rect 119246 124584 119252 124636
rect 119304 124624 119310 124636
rect 200298 124624 200304 124636
rect 119304 124596 200304 124624
rect 119304 124584 119310 124596
rect 200298 124584 200304 124596
rect 200356 124584 200362 124636
rect 121270 124516 121276 124568
rect 121328 124556 121334 124568
rect 202874 124556 202880 124568
rect 121328 124528 202880 124556
rect 121328 124516 121334 124528
rect 202874 124516 202880 124528
rect 202932 124516 202938 124568
rect 119706 124448 119712 124500
rect 119764 124488 119770 124500
rect 201678 124488 201684 124500
rect 119764 124460 201684 124488
rect 119764 124448 119770 124460
rect 201678 124448 201684 124460
rect 201736 124448 201742 124500
rect 115290 124380 115296 124432
rect 115348 124420 115354 124432
rect 203150 124420 203156 124432
rect 115348 124392 203156 124420
rect 115348 124380 115354 124392
rect 203150 124380 203156 124392
rect 203208 124380 203214 124432
rect 108574 124312 108580 124364
rect 108632 124352 108638 124364
rect 201862 124352 201868 124364
rect 108632 124324 201868 124352
rect 108632 124312 108638 124324
rect 201862 124312 201868 124324
rect 201920 124312 201926 124364
rect 108666 124244 108672 124296
rect 108724 124284 108730 124296
rect 203058 124284 203064 124296
rect 108724 124256 203064 124284
rect 108724 124244 108730 124256
rect 203058 124244 203064 124256
rect 203116 124244 203122 124296
rect 174538 124176 174544 124228
rect 174596 124216 174602 124228
rect 306374 124216 306380 124228
rect 174596 124188 306380 124216
rect 174596 124176 174602 124188
rect 306374 124176 306380 124188
rect 306432 124176 306438 124228
rect 109770 124108 109776 124160
rect 109828 124148 109834 124160
rect 110230 124148 110236 124160
rect 109828 124120 110236 124148
rect 109828 124108 109834 124120
rect 110230 124108 110236 124120
rect 110288 124108 110294 124160
rect 119154 124108 119160 124160
rect 119212 124148 119218 124160
rect 119522 124148 119528 124160
rect 119212 124120 119528 124148
rect 119212 124108 119218 124120
rect 119522 124108 119528 124120
rect 119580 124108 119586 124160
rect 120902 124108 120908 124160
rect 120960 124148 120966 124160
rect 121178 124148 121184 124160
rect 120960 124120 121184 124148
rect 120960 124108 120966 124120
rect 121178 124108 121184 124120
rect 121236 124108 121242 124160
rect 164970 124108 164976 124160
rect 165028 124148 165034 124160
rect 165522 124148 165528 124160
rect 165028 124120 165528 124148
rect 165028 124108 165034 124120
rect 165522 124108 165528 124120
rect 165580 124108 165586 124160
rect 182910 124108 182916 124160
rect 182968 124148 182974 124160
rect 183554 124148 183560 124160
rect 182968 124120 183560 124148
rect 182968 124108 182974 124120
rect 183554 124108 183560 124120
rect 183612 124108 183618 124160
rect 202138 124108 202144 124160
rect 202196 124148 202202 124160
rect 202414 124148 202420 124160
rect 202196 124120 202420 124148
rect 202196 124108 202202 124120
rect 202414 124108 202420 124120
rect 202472 124108 202478 124160
rect 208394 124108 208400 124160
rect 208452 124148 208458 124160
rect 209038 124148 209044 124160
rect 208452 124120 209044 124148
rect 208452 124108 208458 124120
rect 209038 124108 209044 124120
rect 209096 124108 209102 124160
rect 167270 123700 167276 123752
rect 167328 123740 167334 123752
rect 167822 123740 167828 123752
rect 167328 123712 167828 123740
rect 167328 123700 167334 123712
rect 167822 123700 167828 123712
rect 167880 123700 167886 123752
rect 165246 123632 165252 123684
rect 165304 123672 165310 123684
rect 201954 123672 201960 123684
rect 165304 123644 201960 123672
rect 165304 123632 165310 123644
rect 201954 123632 201960 123644
rect 202012 123672 202018 123684
rect 229646 123672 229652 123684
rect 202012 123644 229652 123672
rect 202012 123632 202018 123644
rect 229646 123632 229652 123644
rect 229704 123632 229710 123684
rect 165154 123564 165160 123616
rect 165212 123604 165218 123616
rect 202414 123604 202420 123616
rect 165212 123576 202420 123604
rect 165212 123564 165218 123576
rect 202414 123564 202420 123576
rect 202472 123564 202478 123616
rect 165062 123496 165068 123548
rect 165120 123536 165126 123548
rect 202322 123536 202328 123548
rect 165120 123508 202328 123536
rect 165120 123496 165126 123508
rect 202322 123496 202328 123508
rect 202380 123496 202386 123548
rect 3418 123428 3424 123480
rect 3476 123468 3482 123480
rect 95878 123468 95884 123480
rect 3476 123440 95884 123468
rect 3476 123428 3482 123440
rect 95878 123428 95884 123440
rect 95936 123428 95942 123480
rect 112530 123428 112536 123480
rect 112588 123468 112594 123480
rect 112898 123468 112904 123480
rect 112588 123440 112904 123468
rect 112588 123428 112594 123440
rect 112898 123428 112904 123440
rect 112956 123468 112962 123480
rect 229094 123468 229100 123480
rect 112956 123440 229100 123468
rect 112956 123428 112962 123440
rect 229094 123428 229100 123440
rect 229152 123468 229158 123480
rect 229738 123468 229744 123480
rect 229152 123440 229744 123468
rect 229152 123428 229158 123440
rect 229738 123428 229744 123440
rect 229796 123428 229802 123480
rect 159542 123360 159548 123412
rect 159600 123400 159606 123412
rect 205726 123400 205732 123412
rect 159600 123372 205732 123400
rect 159600 123360 159606 123372
rect 205726 123360 205732 123372
rect 205784 123360 205790 123412
rect 162394 123292 162400 123344
rect 162452 123332 162458 123344
rect 208394 123332 208400 123344
rect 162452 123304 208400 123332
rect 162452 123292 162458 123304
rect 208394 123292 208400 123304
rect 208452 123292 208458 123344
rect 119522 123224 119528 123276
rect 119580 123264 119586 123276
rect 200206 123264 200212 123276
rect 119580 123236 200212 123264
rect 119580 123224 119586 123236
rect 200206 123224 200212 123236
rect 200264 123224 200270 123276
rect 120902 123156 120908 123208
rect 120960 123196 120966 123208
rect 204622 123196 204628 123208
rect 120960 123168 204628 123196
rect 120960 123156 120966 123168
rect 204622 123156 204628 123168
rect 204680 123156 204686 123208
rect 119430 123088 119436 123140
rect 119488 123128 119494 123140
rect 119488 123100 122834 123128
rect 119488 123088 119494 123100
rect 122806 123060 122834 123100
rect 164970 123088 164976 123140
rect 165028 123128 165034 123140
rect 175826 123128 175832 123140
rect 165028 123100 175832 123128
rect 165028 123088 165034 123100
rect 175826 123088 175832 123100
rect 175884 123128 175890 123140
rect 259454 123128 259460 123140
rect 175884 123100 259460 123128
rect 175884 123088 175890 123100
rect 259454 123088 259460 123100
rect 259512 123088 259518 123140
rect 204530 123060 204536 123072
rect 122806 123032 204536 123060
rect 204530 123020 204536 123032
rect 204588 123020 204594 123072
rect 115750 122952 115756 123004
rect 115808 122992 115814 123004
rect 204714 122992 204720 123004
rect 115808 122964 204720 122992
rect 115808 122952 115814 122964
rect 204714 122952 204720 122964
rect 204772 122952 204778 123004
rect 112990 122884 112996 122936
rect 113048 122924 113054 122936
rect 203242 122924 203248 122936
rect 113048 122896 203248 122924
rect 113048 122884 113054 122896
rect 203242 122884 203248 122896
rect 203300 122884 203306 122936
rect 109770 122816 109776 122868
rect 109828 122856 109834 122868
rect 202966 122856 202972 122868
rect 109828 122828 112484 122856
rect 109828 122816 109834 122828
rect 112456 122788 112484 122828
rect 113008 122828 202972 122856
rect 113008 122788 113036 122828
rect 202966 122816 202972 122828
rect 203024 122816 203030 122868
rect 112456 122760 113036 122788
rect 170950 122612 170956 122664
rect 171008 122652 171014 122664
rect 197722 122652 197728 122664
rect 171008 122624 197728 122652
rect 171008 122612 171014 122624
rect 197722 122612 197728 122624
rect 197780 122612 197786 122664
rect 179690 122544 179696 122596
rect 179748 122584 179754 122596
rect 187694 122584 187700 122596
rect 179748 122556 187700 122584
rect 179748 122544 179754 122556
rect 187694 122544 187700 122556
rect 187752 122544 187758 122596
rect 155218 122476 155224 122528
rect 155276 122516 155282 122528
rect 187418 122516 187424 122528
rect 155276 122488 187424 122516
rect 155276 122476 155282 122488
rect 187418 122476 187424 122488
rect 187476 122476 187482 122528
rect 88334 122408 88340 122460
rect 88392 122448 88398 122460
rect 131942 122448 131948 122460
rect 88392 122420 131948 122448
rect 88392 122408 88398 122420
rect 131942 122408 131948 122420
rect 132000 122448 132006 122460
rect 181806 122448 181812 122460
rect 132000 122420 181812 122448
rect 132000 122408 132006 122420
rect 181806 122408 181812 122420
rect 181864 122408 181870 122460
rect 92198 122340 92204 122392
rect 92256 122380 92262 122392
rect 130562 122380 130568 122392
rect 92256 122352 130568 122380
rect 92256 122340 92262 122352
rect 130562 122340 130568 122352
rect 130620 122380 130626 122392
rect 184750 122380 184756 122392
rect 130620 122352 184756 122380
rect 130620 122340 130626 122352
rect 184750 122340 184756 122352
rect 184808 122340 184814 122392
rect 99282 122272 99288 122324
rect 99340 122312 99346 122324
rect 159358 122312 159364 122324
rect 99340 122284 159364 122312
rect 99340 122272 99346 122284
rect 159358 122272 159364 122284
rect 159416 122312 159422 122324
rect 159416 122284 161474 122312
rect 159416 122272 159422 122284
rect 93854 122204 93860 122256
rect 93912 122244 93918 122256
rect 155218 122244 155224 122256
rect 93912 122216 155224 122244
rect 93912 122204 93918 122216
rect 155218 122204 155224 122216
rect 155276 122204 155282 122256
rect 161446 122244 161474 122284
rect 163682 122272 163688 122324
rect 163740 122312 163746 122324
rect 164142 122312 164148 122324
rect 163740 122284 164148 122312
rect 163740 122272 163746 122284
rect 164142 122272 164148 122284
rect 164200 122272 164206 122324
rect 173250 122272 173256 122324
rect 173308 122312 173314 122324
rect 292574 122312 292580 122324
rect 173308 122284 292580 122312
rect 173308 122272 173314 122284
rect 292574 122272 292580 122284
rect 292632 122272 292638 122324
rect 191926 122244 191932 122256
rect 161446 122216 191932 122244
rect 191926 122204 191932 122216
rect 191984 122244 191990 122256
rect 325694 122244 325700 122256
rect 191984 122216 325700 122244
rect 191984 122204 191990 122216
rect 325694 122204 325700 122216
rect 325752 122204 325758 122256
rect 91094 122136 91100 122188
rect 91152 122176 91158 122188
rect 159450 122176 159456 122188
rect 91152 122148 159456 122176
rect 91152 122136 91158 122148
rect 159450 122136 159456 122148
rect 159508 122176 159514 122188
rect 185486 122176 185492 122188
rect 159508 122148 185492 122176
rect 159508 122136 159514 122148
rect 185486 122136 185492 122148
rect 185544 122136 185550 122188
rect 188062 122136 188068 122188
rect 188120 122176 188126 122188
rect 198826 122176 198832 122188
rect 188120 122148 198832 122176
rect 188120 122136 188126 122148
rect 198826 122136 198832 122148
rect 198884 122136 198890 122188
rect 117130 122068 117136 122120
rect 117188 122108 117194 122120
rect 226334 122108 226340 122120
rect 117188 122080 226340 122108
rect 117188 122068 117194 122080
rect 226334 122068 226340 122080
rect 226392 122068 226398 122120
rect 166810 122000 166816 122052
rect 166868 122040 166874 122052
rect 193858 122040 193864 122052
rect 166868 122012 193864 122040
rect 166868 122000 166874 122012
rect 193858 122000 193864 122012
rect 193916 122000 193922 122052
rect 184750 121932 184756 121984
rect 184808 121972 184814 121984
rect 200942 121972 200948 121984
rect 184808 121944 200948 121972
rect 184808 121932 184814 121944
rect 200942 121932 200948 121944
rect 201000 121932 201006 121984
rect 187418 121864 187424 121916
rect 187476 121904 187482 121916
rect 203702 121904 203708 121916
rect 187476 121876 203708 121904
rect 187476 121864 187482 121876
rect 203702 121864 203708 121876
rect 203760 121864 203766 121916
rect 181806 121796 181812 121848
rect 181864 121836 181870 121848
rect 200758 121836 200764 121848
rect 181864 121808 200764 121836
rect 181864 121796 181870 121808
rect 200758 121796 200764 121808
rect 200816 121796 200822 121848
rect 163682 121728 163688 121780
rect 163740 121768 163746 121780
rect 175274 121768 175280 121780
rect 163740 121740 175280 121768
rect 163740 121728 163746 121740
rect 175274 121728 175280 121740
rect 175332 121728 175338 121780
rect 186130 121768 186136 121780
rect 180766 121740 186136 121768
rect 169754 121660 169760 121712
rect 169812 121700 169818 121712
rect 180766 121700 180794 121740
rect 186130 121728 186136 121740
rect 186188 121768 186194 121780
rect 186188 121740 195284 121768
rect 186188 121728 186194 121740
rect 169812 121672 180794 121700
rect 169812 121660 169818 121672
rect 184842 121660 184848 121712
rect 184900 121700 184906 121712
rect 190638 121700 190644 121712
rect 184900 121672 190644 121700
rect 184900 121660 184906 121672
rect 190638 121660 190644 121672
rect 190696 121660 190702 121712
rect 195256 121700 195284 121740
rect 196434 121728 196440 121780
rect 196492 121768 196498 121780
rect 206278 121768 206284 121780
rect 196492 121740 206284 121768
rect 196492 121728 196498 121740
rect 206278 121728 206284 121740
rect 206336 121728 206342 121780
rect 220078 121700 220084 121712
rect 195256 121672 220084 121700
rect 220078 121660 220084 121672
rect 220136 121660 220142 121712
rect 226334 121660 226340 121712
rect 226392 121700 226398 121712
rect 226978 121700 226984 121712
rect 226392 121672 226984 121700
rect 226392 121660 226398 121672
rect 226978 121660 226984 121672
rect 227036 121660 227042 121712
rect 104894 121592 104900 121644
rect 104952 121632 104958 121644
rect 199010 121632 199016 121644
rect 104952 121604 199016 121632
rect 104952 121592 104958 121604
rect 199010 121592 199016 121604
rect 199068 121632 199074 121644
rect 199838 121632 199844 121644
rect 199068 121604 199844 121632
rect 199068 121592 199074 121604
rect 199838 121592 199844 121604
rect 199896 121632 199902 121644
rect 313274 121632 313280 121644
rect 199896 121604 313280 121632
rect 199896 121592 199902 121604
rect 313274 121592 313280 121604
rect 313332 121592 313338 121644
rect 186222 121524 186228 121576
rect 186280 121564 186286 121576
rect 188062 121564 188068 121576
rect 186280 121536 188068 121564
rect 186280 121524 186286 121536
rect 188062 121524 188068 121536
rect 188120 121524 188126 121576
rect 196434 121564 196440 121576
rect 190426 121536 196440 121564
rect 116762 121456 116768 121508
rect 116820 121496 116826 121508
rect 117130 121496 117136 121508
rect 116820 121468 117136 121496
rect 116820 121456 116826 121468
rect 117130 121456 117136 121468
rect 117188 121456 117194 121508
rect 169846 121456 169852 121508
rect 169904 121496 169910 121508
rect 183554 121496 183560 121508
rect 169904 121468 183560 121496
rect 169904 121456 169910 121468
rect 183554 121456 183560 121468
rect 183612 121456 183618 121508
rect 186314 121456 186320 121508
rect 186372 121496 186378 121508
rect 190426 121496 190454 121536
rect 196434 121524 196440 121536
rect 196492 121524 196498 121576
rect 186372 121468 190454 121496
rect 186372 121456 186378 121468
rect 193122 121456 193128 121508
rect 193180 121496 193186 121508
rect 197078 121496 197084 121508
rect 193180 121468 197084 121496
rect 193180 121456 193186 121468
rect 197078 121456 197084 121468
rect 197136 121456 197142 121508
rect 102410 121388 102416 121440
rect 102468 121428 102474 121440
rect 131114 121428 131120 121440
rect 102468 121400 131120 121428
rect 102468 121388 102474 121400
rect 131114 121388 131120 121400
rect 131172 121388 131178 121440
rect 143442 121388 143448 121440
rect 143500 121428 143506 121440
rect 177114 121428 177120 121440
rect 143500 121400 177120 121428
rect 143500 121388 143506 121400
rect 177114 121388 177120 121400
rect 177172 121388 177178 121440
rect 103790 121320 103796 121372
rect 103848 121360 103854 121372
rect 144178 121360 144184 121372
rect 103848 121332 144184 121360
rect 103848 121320 103854 121332
rect 144178 121320 144184 121332
rect 144236 121320 144242 121372
rect 148318 121320 148324 121372
rect 148376 121360 148382 121372
rect 179690 121360 179696 121372
rect 148376 121332 179696 121360
rect 148376 121320 148382 121332
rect 179690 121320 179696 121332
rect 179748 121320 179754 121372
rect 95418 121252 95424 121304
rect 95476 121292 95482 121304
rect 140038 121292 140044 121304
rect 95476 121264 140044 121292
rect 95476 121252 95482 121264
rect 140038 121252 140044 121264
rect 140096 121292 140102 121304
rect 189994 121292 190000 121304
rect 140096 121264 190000 121292
rect 140096 121252 140102 121264
rect 189994 121252 190000 121264
rect 190052 121252 190058 121304
rect 102134 121184 102140 121236
rect 102192 121224 102198 121236
rect 162118 121224 162124 121236
rect 102192 121196 162124 121224
rect 102192 121184 102198 121196
rect 162118 121184 162124 121196
rect 162176 121224 162182 121236
rect 186314 121224 186320 121236
rect 162176 121196 186320 121224
rect 162176 121184 162182 121196
rect 186314 121184 186320 121196
rect 186372 121184 186378 121236
rect 83090 121116 83096 121168
rect 83148 121156 83154 121168
rect 142890 121156 142896 121168
rect 83148 121128 142896 121156
rect 83148 121116 83154 121128
rect 142890 121116 142896 121128
rect 142948 121156 142954 121168
rect 143442 121156 143448 121168
rect 142948 121128 143448 121156
rect 142948 121116 142954 121128
rect 143442 121116 143448 121128
rect 143500 121116 143506 121168
rect 144178 121116 144184 121168
rect 144236 121156 144242 121168
rect 198366 121156 198372 121168
rect 144236 121128 198372 121156
rect 144236 121116 144242 121128
rect 198366 121116 198372 121128
rect 198424 121116 198430 121168
rect 85574 121048 85580 121100
rect 85632 121088 85638 121100
rect 148318 121088 148324 121100
rect 85632 121060 148324 121088
rect 85632 121048 85638 121060
rect 148318 121048 148324 121060
rect 148376 121048 148382 121100
rect 186222 121088 186228 121100
rect 156616 121060 186228 121088
rect 156616 121032 156644 121060
rect 186222 121048 186228 121060
rect 186280 121048 186286 121100
rect 94130 120980 94136 121032
rect 94188 121020 94194 121032
rect 156598 121020 156604 121032
rect 94188 120992 156604 121020
rect 94188 120980 94194 120992
rect 156598 120980 156604 120992
rect 156656 120980 156662 121032
rect 158070 120980 158076 121032
rect 158128 121020 158134 121032
rect 173250 121020 173256 121032
rect 158128 120992 173256 121020
rect 158128 120980 158134 120992
rect 173250 120980 173256 120992
rect 173308 120980 173314 121032
rect 80514 120912 80520 120964
rect 80572 120952 80578 120964
rect 146938 120952 146944 120964
rect 80572 120924 146944 120952
rect 80572 120912 80578 120924
rect 146938 120912 146944 120924
rect 146996 120952 147002 120964
rect 174538 120952 174544 120964
rect 146996 120924 174544 120952
rect 146996 120912 147002 120924
rect 174538 120912 174544 120924
rect 174596 120912 174602 120964
rect 120718 120844 120724 120896
rect 120776 120884 120782 120896
rect 227714 120884 227720 120896
rect 120776 120856 227720 120884
rect 120776 120844 120782 120856
rect 227714 120844 227720 120856
rect 227772 120844 227778 120896
rect 84194 120776 84200 120828
rect 84252 120816 84258 120828
rect 151078 120816 151084 120828
rect 84252 120788 151084 120816
rect 84252 120776 84258 120788
rect 151078 120776 151084 120788
rect 151136 120816 151142 120828
rect 177758 120816 177764 120828
rect 151136 120788 177764 120816
rect 151136 120776 151142 120788
rect 177758 120776 177764 120788
rect 177816 120816 177822 120828
rect 177816 120788 180794 120816
rect 177816 120776 177822 120788
rect 86862 120708 86868 120760
rect 86920 120748 86926 120760
rect 158070 120748 158076 120760
rect 86920 120720 158076 120748
rect 86920 120708 86926 120720
rect 158070 120708 158076 120720
rect 158128 120708 158134 120760
rect 180766 120748 180794 120788
rect 187694 120776 187700 120828
rect 187752 120816 187758 120828
rect 299474 120816 299480 120828
rect 187752 120788 299480 120816
rect 187752 120776 187758 120788
rect 299474 120776 299480 120788
rect 299532 120776 299538 120828
rect 304994 120748 305000 120760
rect 180766 120720 305000 120748
rect 304994 120708 305000 120720
rect 305052 120708 305058 120760
rect 169754 120640 169760 120692
rect 169812 120680 169818 120692
rect 184842 120680 184848 120692
rect 169812 120652 184848 120680
rect 169812 120640 169818 120652
rect 184842 120640 184848 120652
rect 184900 120640 184906 120692
rect 166166 120572 166172 120624
rect 166224 120612 166230 120624
rect 195146 120612 195152 120624
rect 166224 120584 195152 120612
rect 166224 120572 166230 120584
rect 195146 120572 195152 120584
rect 195204 120572 195210 120624
rect 186774 120504 186780 120556
rect 186832 120544 186838 120556
rect 203610 120544 203616 120556
rect 186832 120516 203616 120544
rect 186832 120504 186838 120516
rect 203610 120504 203616 120516
rect 203668 120504 203674 120556
rect 177114 120436 177120 120488
rect 177172 120476 177178 120488
rect 203518 120476 203524 120488
rect 177172 120448 203524 120476
rect 177172 120436 177178 120448
rect 203518 120436 203524 120448
rect 203576 120436 203582 120488
rect 166074 120368 166080 120420
rect 166132 120408 166138 120420
rect 195054 120408 195060 120420
rect 166132 120380 195060 120408
rect 166132 120368 166138 120380
rect 195054 120368 195060 120380
rect 195112 120408 195118 120420
rect 195790 120408 195796 120420
rect 195112 120380 195796 120408
rect 195112 120368 195118 120380
rect 195790 120368 195796 120380
rect 195848 120368 195854 120420
rect 227714 120368 227720 120420
rect 227772 120408 227778 120420
rect 228726 120408 228732 120420
rect 227772 120380 228732 120408
rect 227772 120368 227778 120380
rect 228726 120368 228732 120380
rect 228784 120368 228790 120420
rect 168558 120300 168564 120352
rect 168616 120340 168622 120352
rect 168616 120312 170076 120340
rect 168616 120300 168622 120312
rect 169938 120272 169944 120284
rect 169496 120244 169944 120272
rect 161446 120040 166396 120068
rect 133230 120000 133236 120012
rect 122806 119972 133236 120000
rect 103606 119688 103612 119740
rect 103664 119728 103670 119740
rect 122806 119728 122834 119972
rect 133230 119960 133236 119972
rect 133288 120000 133294 120012
rect 161446 120000 161474 120040
rect 133288 119972 161474 120000
rect 166368 120000 166396 120040
rect 166442 120028 166448 120080
rect 166500 120068 166506 120080
rect 169496 120068 169524 120244
rect 169938 120232 169944 120244
rect 169996 120232 170002 120284
rect 170048 120204 170076 120312
rect 193858 120300 193864 120352
rect 193916 120340 193922 120352
rect 252554 120340 252560 120352
rect 193916 120312 252560 120340
rect 193916 120300 193922 120312
rect 252554 120300 252560 120312
rect 252612 120300 252618 120352
rect 175274 120232 175280 120284
rect 175332 120272 175338 120284
rect 176470 120272 176476 120284
rect 175332 120244 176476 120272
rect 175332 120232 175338 120244
rect 176470 120232 176476 120244
rect 176528 120272 176534 120284
rect 235258 120272 235264 120284
rect 176528 120244 235264 120272
rect 176528 120232 176534 120244
rect 235258 120232 235264 120244
rect 235316 120232 235322 120284
rect 182910 120204 182916 120216
rect 170048 120176 182916 120204
rect 182910 120164 182916 120176
rect 182968 120164 182974 120216
rect 185486 120164 185492 120216
rect 185544 120204 185550 120216
rect 295334 120204 295340 120216
rect 185544 120176 295340 120204
rect 185544 120164 185550 120176
rect 295334 120164 295340 120176
rect 295392 120164 295398 120216
rect 193214 120096 193220 120148
rect 193272 120136 193278 120148
rect 580350 120136 580356 120148
rect 193272 120108 580356 120136
rect 193272 120096 193278 120108
rect 580350 120096 580356 120108
rect 580408 120096 580414 120148
rect 170950 120068 170956 120080
rect 166500 120040 169524 120068
rect 169772 120040 170956 120068
rect 166500 120028 166506 120040
rect 169772 120000 169800 120040
rect 170950 120028 170956 120040
rect 171008 120028 171014 120080
rect 166368 119972 169800 120000
rect 133288 119960 133294 119972
rect 135162 119892 135168 119944
rect 135220 119932 135226 119944
rect 169754 119932 169760 119944
rect 135220 119904 169760 119932
rect 135220 119892 135226 119904
rect 169754 119892 169760 119904
rect 169812 119892 169818 119944
rect 169846 119892 169852 119944
rect 169904 119932 169910 119944
rect 171962 119932 171968 119944
rect 169904 119904 171968 119932
rect 169904 119892 169910 119904
rect 171962 119892 171968 119904
rect 172020 119892 172026 119944
rect 199654 119892 199660 119944
rect 199712 119932 199718 119944
rect 200574 119932 200580 119944
rect 199712 119904 200580 119932
rect 199712 119892 199718 119904
rect 200574 119892 200580 119904
rect 200632 119892 200638 119944
rect 166442 119864 166448 119876
rect 103664 119700 122834 119728
rect 132466 119836 166448 119864
rect 103664 119688 103670 119700
rect 86954 119620 86960 119672
rect 87012 119660 87018 119672
rect 130470 119660 130476 119672
rect 87012 119632 130476 119660
rect 87012 119620 87018 119632
rect 130470 119620 130476 119632
rect 130528 119660 130534 119672
rect 132466 119660 132494 119836
rect 166442 119824 166448 119836
rect 166500 119824 166506 119876
rect 169110 119824 169116 119876
rect 169168 119864 169174 119876
rect 171042 119864 171048 119876
rect 169168 119836 171048 119864
rect 169168 119824 169174 119836
rect 171042 119824 171048 119836
rect 171100 119824 171106 119876
rect 172422 119824 172428 119876
rect 172480 119824 172486 119876
rect 197814 119824 197820 119876
rect 197872 119864 197878 119876
rect 197872 119836 198780 119864
rect 197872 119824 197878 119836
rect 172440 119796 172468 119824
rect 169772 119768 172468 119796
rect 166626 119688 166632 119740
rect 166684 119728 166690 119740
rect 166902 119728 166908 119740
rect 166684 119700 166908 119728
rect 166684 119688 166690 119700
rect 166902 119688 166908 119700
rect 166960 119728 166966 119740
rect 169662 119728 169668 119740
rect 166960 119700 169668 119728
rect 166960 119688 166966 119700
rect 169662 119688 169668 119700
rect 169720 119688 169726 119740
rect 130528 119632 132494 119660
rect 130528 119620 130534 119632
rect 89714 119552 89720 119604
rect 89772 119592 89778 119604
rect 134610 119592 134616 119604
rect 89772 119564 134616 119592
rect 89772 119552 89778 119564
rect 134610 119552 134616 119564
rect 134668 119592 134674 119604
rect 135162 119592 135168 119604
rect 134668 119564 135168 119592
rect 134668 119552 134674 119564
rect 135162 119552 135168 119564
rect 135220 119552 135226 119604
rect 169772 119592 169800 119768
rect 169846 119688 169852 119740
rect 169904 119688 169910 119740
rect 161446 119564 169800 119592
rect 79318 119484 79324 119536
rect 79376 119524 79382 119536
rect 161446 119524 161474 119564
rect 79376 119496 161474 119524
rect 79376 119484 79382 119496
rect 78490 119416 78496 119468
rect 78548 119456 78554 119468
rect 169864 119456 169892 119688
rect 78548 119428 169892 119456
rect 78548 119416 78554 119428
rect 78582 119348 78588 119400
rect 78640 119388 78646 119400
rect 169110 119388 169116 119400
rect 78640 119360 169116 119388
rect 78640 119348 78646 119360
rect 169110 119348 169116 119360
rect 169168 119348 169174 119400
rect 198752 119388 198780 119836
rect 198826 119824 198832 119876
rect 198884 119864 198890 119876
rect 198884 119836 200114 119864
rect 198884 119824 198890 119836
rect 200086 119456 200114 119836
rect 251174 119456 251180 119468
rect 200086 119428 251180 119456
rect 251174 119416 251180 119428
rect 251232 119416 251238 119468
rect 271874 119388 271880 119400
rect 198752 119360 271880 119388
rect 271874 119348 271880 119360
rect 271932 119348 271938 119400
rect 167270 119280 167276 119332
rect 167328 119320 167334 119332
rect 169662 119320 169668 119332
rect 167328 119292 169668 119320
rect 167328 119280 167334 119292
rect 169662 119280 169668 119292
rect 169720 119280 169726 119332
rect 200574 118980 200580 118992
rect 180766 118952 200580 118980
rect 166442 118872 166448 118924
rect 166500 118912 166506 118924
rect 180766 118912 180794 118952
rect 200574 118940 200580 118952
rect 200632 118940 200638 118992
rect 166500 118884 180794 118912
rect 166500 118872 166506 118884
rect 165338 118804 165344 118856
rect 165396 118844 165402 118856
rect 200114 118844 200120 118856
rect 165396 118816 200120 118844
rect 165396 118804 165402 118816
rect 200086 118804 200120 118816
rect 200172 118804 200178 118856
rect 200086 118708 200114 118804
rect 349154 118708 349160 118720
rect 200086 118680 349160 118708
rect 349154 118668 349160 118680
rect 349212 118668 349218 118720
rect 64690 118600 64696 118652
rect 64748 118640 64754 118652
rect 78490 118640 78496 118652
rect 64748 118612 78496 118640
rect 64748 118600 64754 118612
rect 78490 118600 78496 118612
rect 78548 118600 78554 118652
rect 138106 118600 138112 118652
rect 138164 118640 138170 118652
rect 138658 118640 138664 118652
rect 138164 118612 138664 118640
rect 138164 118600 138170 118612
rect 138658 118600 138664 118612
rect 138716 118640 138722 118652
rect 164142 118640 164148 118652
rect 138716 118612 164148 118640
rect 138716 118600 138722 118612
rect 164142 118600 164148 118612
rect 164200 118600 164206 118652
rect 167178 118600 167184 118652
rect 167236 118640 167242 118652
rect 167730 118640 167736 118652
rect 167236 118612 167736 118640
rect 167236 118600 167242 118612
rect 167730 118600 167736 118612
rect 167788 118600 167794 118652
rect 65978 118532 65984 118584
rect 66036 118572 66042 118584
rect 77754 118572 77760 118584
rect 66036 118544 77760 118572
rect 66036 118532 66042 118544
rect 77754 118532 77760 118544
rect 77812 118572 77818 118584
rect 78582 118572 78588 118584
rect 77812 118544 78588 118572
rect 77812 118532 77818 118544
rect 78582 118532 78588 118544
rect 78640 118532 78646 118584
rect 157334 118532 157340 118584
rect 157392 118572 157398 118584
rect 157978 118572 157984 118584
rect 157392 118544 157984 118572
rect 157392 118532 157398 118544
rect 157978 118532 157984 118544
rect 158036 118572 158042 118584
rect 169754 118572 169760 118584
rect 158036 118544 169760 118572
rect 158036 118532 158042 118544
rect 169754 118532 169760 118544
rect 169812 118532 169818 118584
rect 92474 118056 92480 118108
rect 92532 118096 92538 118108
rect 138106 118096 138112 118108
rect 92532 118068 138112 118096
rect 92532 118056 92538 118068
rect 138106 118056 138112 118068
rect 138164 118056 138170 118108
rect 164786 118056 164792 118108
rect 164844 118096 164850 118108
rect 165154 118096 165160 118108
rect 164844 118068 165160 118096
rect 164844 118056 164850 118068
rect 165154 118056 165160 118068
rect 165212 118056 165218 118108
rect 91554 117988 91560 118040
rect 91612 118028 91618 118040
rect 157334 118028 157340 118040
rect 91612 118000 157340 118028
rect 91612 117988 91618 118000
rect 157334 117988 157340 118000
rect 157392 117988 157398 118040
rect 99834 117920 99840 117972
rect 99892 117960 99898 117972
rect 166810 117960 166816 117972
rect 99892 117932 166816 117960
rect 99892 117920 99898 117932
rect 166810 117920 166816 117932
rect 166868 117920 166874 117972
rect 201954 117920 201960 117972
rect 202012 117960 202018 117972
rect 202874 117960 202880 117972
rect 202012 117932 202880 117960
rect 202012 117920 202018 117932
rect 202874 117920 202880 117932
rect 202932 117960 202938 117972
rect 580258 117960 580264 117972
rect 202932 117932 580264 117960
rect 202932 117920 202938 117932
rect 580258 117920 580264 117932
rect 580316 117920 580322 117972
rect 80054 117444 80060 117496
rect 80112 117484 80118 117496
rect 167086 117484 167092 117496
rect 80112 117456 167092 117484
rect 80112 117444 80118 117456
rect 167086 117444 167092 117456
rect 167144 117444 167150 117496
rect 75914 117376 75920 117428
rect 75972 117416 75978 117428
rect 166994 117416 167000 117428
rect 75972 117388 167000 117416
rect 75972 117376 75978 117388
rect 166994 117376 167000 117388
rect 167052 117376 167058 117428
rect 65978 117308 65984 117360
rect 66036 117348 66042 117360
rect 167914 117348 167920 117360
rect 66036 117320 167920 117348
rect 66036 117308 66042 117320
rect 167914 117308 167920 117320
rect 167972 117308 167978 117360
rect 63310 117240 63316 117292
rect 63368 117280 63374 117292
rect 76466 117280 76472 117292
rect 63368 117252 76472 117280
rect 63368 117240 63374 117252
rect 76466 117240 76472 117252
rect 76524 117280 76530 117292
rect 77110 117280 77116 117292
rect 76524 117252 77116 117280
rect 76524 117240 76530 117252
rect 77110 117240 77116 117252
rect 77168 117240 77174 117292
rect 126238 117240 126244 117292
rect 126296 117280 126302 117292
rect 126790 117280 126796 117292
rect 126296 117252 126796 117280
rect 126296 117240 126302 117252
rect 126790 117240 126796 117252
rect 126848 117280 126854 117292
rect 166534 117280 166540 117292
rect 126848 117252 166540 117280
rect 126848 117240 126854 117252
rect 166534 117240 166540 117252
rect 166592 117240 166598 117292
rect 64782 117172 64788 117224
rect 64840 117212 64846 117224
rect 75914 117212 75920 117224
rect 64840 117184 75920 117212
rect 64840 117172 64846 117184
rect 75914 117172 75920 117184
rect 75972 117172 75978 117224
rect 137370 117172 137376 117224
rect 137428 117212 137434 117224
rect 168650 117212 168656 117224
rect 137428 117184 168656 117212
rect 137428 117172 137434 117184
rect 168650 117172 168656 117184
rect 168708 117172 168714 117224
rect 97994 116696 98000 116748
rect 98052 116736 98058 116748
rect 137370 116736 137376 116748
rect 98052 116708 137376 116736
rect 98052 116696 98058 116708
rect 137370 116696 137376 116708
rect 137428 116696 137434 116748
rect 84378 116628 84384 116680
rect 84436 116668 84442 116680
rect 126790 116668 126796 116680
rect 84436 116640 126796 116668
rect 84436 116628 84442 116640
rect 126790 116628 126796 116640
rect 126848 116628 126854 116680
rect 82906 116560 82912 116612
rect 82964 116600 82970 116612
rect 163682 116600 163688 116612
rect 82964 116572 163688 116600
rect 82964 116560 82970 116572
rect 163682 116560 163688 116572
rect 163740 116560 163746 116612
rect 202138 116560 202144 116612
rect 202196 116600 202202 116612
rect 202966 116600 202972 116612
rect 202196 116572 202972 116600
rect 202196 116560 202202 116572
rect 202966 116560 202972 116572
rect 203024 116600 203030 116612
rect 282914 116600 282920 116612
rect 203024 116572 282920 116600
rect 203024 116560 203030 116572
rect 282914 116560 282920 116572
rect 282972 116560 282978 116612
rect 72602 116084 72608 116136
rect 72660 116124 72666 116136
rect 169110 116124 169116 116136
rect 72660 116096 169116 116124
rect 72660 116084 72666 116096
rect 169110 116084 169116 116096
rect 169168 116084 169174 116136
rect 64414 116016 64420 116068
rect 64472 116056 64478 116068
rect 167638 116056 167644 116068
rect 64472 116028 167644 116056
rect 64472 116016 64478 116028
rect 167638 116016 167644 116028
rect 167696 116016 167702 116068
rect 64690 115948 64696 116000
rect 64748 115988 64754 116000
rect 167730 115988 167736 116000
rect 64748 115960 167736 115988
rect 64748 115948 64754 115960
rect 167730 115948 167736 115960
rect 167788 115948 167794 116000
rect 97718 115880 97724 115932
rect 97776 115920 97782 115932
rect 99282 115920 99288 115932
rect 97776 115892 99288 115920
rect 97776 115880 97782 115892
rect 99282 115880 99288 115892
rect 99340 115880 99346 115932
rect 134610 115880 134616 115932
rect 134668 115920 134674 115932
rect 165982 115920 165988 115932
rect 134668 115892 165988 115920
rect 134668 115880 134674 115892
rect 165982 115880 165988 115892
rect 166040 115880 166046 115932
rect 144914 115812 144920 115864
rect 144972 115852 144978 115864
rect 145558 115852 145564 115864
rect 144972 115824 145564 115852
rect 144972 115812 144978 115824
rect 145558 115812 145564 115824
rect 145616 115812 145622 115864
rect 154574 115608 154580 115660
rect 154632 115648 154638 115660
rect 155218 115648 155224 115660
rect 154632 115620 155224 115648
rect 154632 115608 154638 115620
rect 155218 115608 155224 115620
rect 155276 115608 155282 115660
rect 97074 115336 97080 115388
rect 97132 115376 97138 115388
rect 134610 115376 134616 115388
rect 97132 115348 134616 115376
rect 97132 115336 97138 115348
rect 134610 115336 134616 115348
rect 134668 115336 134674 115388
rect 75546 115268 75552 115320
rect 75604 115308 75610 115320
rect 80054 115308 80060 115320
rect 75604 115280 80060 115308
rect 75604 115268 75610 115280
rect 80054 115268 80060 115280
rect 80112 115268 80118 115320
rect 82262 115268 82268 115320
rect 82320 115308 82326 115320
rect 164970 115308 164976 115320
rect 82320 115280 164976 115308
rect 82320 115268 82326 115280
rect 164970 115268 164976 115280
rect 165028 115268 165034 115320
rect 75822 115200 75828 115252
rect 75880 115240 75886 115252
rect 166902 115240 166908 115252
rect 75880 115212 166908 115240
rect 75880 115200 75886 115212
rect 166902 115200 166908 115212
rect 166960 115200 166966 115252
rect 201954 115200 201960 115252
rect 202012 115240 202018 115252
rect 203242 115240 203248 115252
rect 202012 115212 203248 115240
rect 202012 115200 202018 115212
rect 203242 115200 203248 115212
rect 203300 115240 203306 115252
rect 314654 115240 314660 115252
rect 203300 115212 314660 115240
rect 203300 115200 203306 115212
rect 314654 115200 314660 115212
rect 314712 115200 314718 115252
rect 64322 115064 64328 115116
rect 64380 115104 64386 115116
rect 145558 115104 145564 115116
rect 64380 115076 145564 115104
rect 64380 115064 64386 115076
rect 145558 115064 145564 115076
rect 145616 115064 145622 115116
rect 69566 114996 69572 115048
rect 69624 115036 69630 115048
rect 154574 115036 154580 115048
rect 69624 115008 154580 115036
rect 69624 114996 69630 115008
rect 154574 114996 154580 115008
rect 154632 114996 154638 115048
rect 73062 114928 73068 114980
rect 73120 114968 73126 114980
rect 166994 114968 167000 114980
rect 73120 114940 167000 114968
rect 73120 114928 73126 114940
rect 166994 114928 167000 114940
rect 167052 114928 167058 114980
rect 71682 114860 71688 114912
rect 71740 114900 71746 114912
rect 167178 114900 167184 114912
rect 71740 114872 167184 114900
rect 71740 114860 71746 114872
rect 167178 114860 167184 114872
rect 167236 114860 167242 114912
rect 66162 114792 66168 114844
rect 66220 114832 66226 114844
rect 162854 114832 162860 114844
rect 66220 114804 162860 114832
rect 66220 114792 66226 114804
rect 162854 114792 162860 114804
rect 162912 114832 162918 114844
rect 163498 114832 163504 114844
rect 162912 114804 163504 114832
rect 162912 114792 162918 114804
rect 163498 114792 163504 114804
rect 163556 114792 163562 114844
rect 64230 114724 64236 114776
rect 64288 114764 64294 114776
rect 162302 114764 162308 114776
rect 64288 114736 162308 114764
rect 64288 114724 64294 114736
rect 162302 114724 162308 114736
rect 162360 114764 162366 114776
rect 162670 114764 162676 114776
rect 162360 114736 162676 114764
rect 162360 114724 162366 114736
rect 162670 114724 162676 114736
rect 162728 114724 162734 114776
rect 70210 114656 70216 114708
rect 70268 114696 70274 114708
rect 167086 114696 167092 114708
rect 70268 114668 167092 114696
rect 70268 114656 70274 114668
rect 167086 114656 167092 114668
rect 167144 114656 167150 114708
rect 65702 114588 65708 114640
rect 65760 114628 65766 114640
rect 167822 114628 167828 114640
rect 65760 114600 167828 114628
rect 65760 114588 65766 114600
rect 167822 114588 167828 114600
rect 167880 114588 167886 114640
rect 64782 114520 64788 114572
rect 64840 114560 64846 114572
rect 167546 114560 167552 114572
rect 64840 114532 167552 114560
rect 64840 114520 64846 114532
rect 167546 114520 167552 114532
rect 167604 114520 167610 114572
rect 60734 114452 60740 114504
rect 60792 114492 60798 114504
rect 62022 114492 62028 114504
rect 60792 114464 62028 114492
rect 60792 114452 60798 114464
rect 62022 114452 62028 114464
rect 62080 114492 62086 114504
rect 79318 114492 79324 114504
rect 62080 114464 79324 114492
rect 62080 114452 62086 114464
rect 79318 114452 79324 114464
rect 79376 114452 79382 114504
rect 95878 114452 95884 114504
rect 95936 114492 95942 114504
rect 96430 114492 96436 114504
rect 95936 114464 96436 114492
rect 95936 114452 95942 114464
rect 96430 114452 96436 114464
rect 96488 114492 96494 114504
rect 124306 114492 124312 114504
rect 96488 114464 124312 114492
rect 96488 114452 96494 114464
rect 124306 114452 124312 114464
rect 124364 114492 124370 114504
rect 166626 114492 166632 114504
rect 124364 114464 166632 114492
rect 124364 114452 124370 114464
rect 166626 114452 166632 114464
rect 166684 114452 166690 114504
rect 65518 114384 65524 114436
rect 65576 114424 65582 114436
rect 75822 114424 75828 114436
rect 65576 114396 75828 114424
rect 65576 114384 65582 114396
rect 75822 114384 75828 114396
rect 75880 114384 75886 114436
rect 90634 114384 90640 114436
rect 90692 114424 90698 114436
rect 92198 114424 92204 114436
rect 90692 114396 92204 114424
rect 90692 114384 90698 114396
rect 92198 114384 92204 114396
rect 92256 114384 92262 114436
rect 124214 114424 124220 114436
rect 122806 114396 124220 114424
rect 61930 114316 61936 114368
rect 61988 114356 61994 114368
rect 71314 114356 71320 114368
rect 61988 114328 71320 114356
rect 61988 114316 61994 114328
rect 71314 114316 71320 114328
rect 71372 114356 71378 114368
rect 71682 114356 71688 114368
rect 71372 114328 71688 114356
rect 71372 114316 71378 114328
rect 71682 114316 71688 114328
rect 71740 114316 71746 114368
rect 74534 114316 74540 114368
rect 74592 114356 74598 114368
rect 75914 114356 75920 114368
rect 74592 114328 75920 114356
rect 74592 114316 74598 114328
rect 75914 114316 75920 114328
rect 75972 114316 75978 114368
rect 67266 114248 67272 114300
rect 67324 114288 67330 114300
rect 67542 114288 67548 114300
rect 67324 114260 67548 114288
rect 67324 114248 67330 114260
rect 67542 114248 67548 114260
rect 67600 114248 67606 114300
rect 100938 114248 100944 114300
rect 100996 114288 101002 114300
rect 122806 114288 122834 114396
rect 124214 114384 124220 114396
rect 124272 114424 124278 114436
rect 166166 114424 166172 114436
rect 124272 114396 166172 114424
rect 124272 114384 124278 114396
rect 166166 114384 166172 114396
rect 166224 114384 166230 114436
rect 127618 114316 127624 114368
rect 127676 114356 127682 114368
rect 168466 114356 168472 114368
rect 127676 114328 168472 114356
rect 127676 114316 127682 114328
rect 168466 114316 168472 114328
rect 168524 114316 168530 114368
rect 126974 114288 126980 114300
rect 100996 114260 122834 114288
rect 123496 114260 126980 114288
rect 100996 114248 101002 114260
rect 66070 114180 66076 114232
rect 66128 114220 66134 114232
rect 71958 114220 71964 114232
rect 66128 114192 71964 114220
rect 66128 114180 66134 114192
rect 71958 114180 71964 114192
rect 72016 114220 72022 114232
rect 73062 114220 73068 114232
rect 72016 114192 73068 114220
rect 72016 114180 72022 114192
rect 73062 114180 73068 114192
rect 73120 114180 73126 114232
rect 101582 114180 101588 114232
rect 101640 114220 101646 114232
rect 123496 114220 123524 114260
rect 126974 114248 126980 114260
rect 127032 114288 127038 114300
rect 166074 114288 166080 114300
rect 127032 114260 166080 114288
rect 127032 114248 127038 114260
rect 166074 114248 166080 114260
rect 166132 114248 166138 114300
rect 133138 114220 133144 114232
rect 101640 114192 123524 114220
rect 132466 114192 133144 114220
rect 101640 114180 101646 114192
rect 95142 114112 95148 114164
rect 95200 114152 95206 114164
rect 132466 114152 132494 114192
rect 133138 114180 133144 114192
rect 133196 114220 133202 114232
rect 168374 114220 168380 114232
rect 133196 114192 168380 114220
rect 133196 114180 133202 114192
rect 168374 114180 168380 114192
rect 168432 114180 168438 114232
rect 95200 114124 132494 114152
rect 95200 114112 95206 114124
rect 86126 114044 86132 114096
rect 86184 114084 86190 114096
rect 127618 114084 127624 114096
rect 86184 114056 127624 114084
rect 86184 114044 86190 114056
rect 127618 114044 127624 114056
rect 127676 114044 127682 114096
rect 99006 113976 99012 114028
rect 99064 114016 99070 114028
rect 142798 114016 142804 114028
rect 99064 113988 142804 114016
rect 99064 113976 99070 113988
rect 142798 113976 142804 113988
rect 142856 114016 142862 114028
rect 143442 114016 143448 114028
rect 142856 113988 143448 114016
rect 142856 113976 142862 113988
rect 143442 113976 143448 113988
rect 143500 113976 143506 114028
rect 81618 113908 81624 113960
rect 81676 113948 81682 113960
rect 140774 113948 140780 113960
rect 81676 113920 140780 113948
rect 81676 113908 81682 113920
rect 140774 113908 140780 113920
rect 140832 113908 140838 113960
rect 88702 113840 88708 113892
rect 88760 113880 88766 113892
rect 152458 113880 152464 113892
rect 88760 113852 152464 113880
rect 88760 113840 88766 113852
rect 152458 113840 152464 113852
rect 152516 113880 152522 113892
rect 153010 113880 153016 113892
rect 152516 113852 153016 113880
rect 152516 113840 152522 113852
rect 153010 113840 153016 113852
rect 153068 113840 153074 113892
rect 3510 113772 3516 113824
rect 3568 113812 3574 113824
rect 60734 113812 60740 113824
rect 3568 113784 60740 113812
rect 3568 113772 3574 113784
rect 60734 113772 60740 113784
rect 60792 113772 60798 113824
rect 64598 113772 64604 113824
rect 64656 113812 64662 113824
rect 69382 113812 69388 113824
rect 64656 113784 69388 113812
rect 64656 113772 64662 113784
rect 69382 113772 69388 113784
rect 69440 113772 69446 113824
rect 89346 113772 89352 113824
rect 89404 113812 89410 113824
rect 168558 113812 168564 113824
rect 89404 113784 168564 113812
rect 89404 113772 89410 113784
rect 168558 113772 168564 113784
rect 168616 113772 168622 113824
rect 200942 113772 200948 113824
rect 201000 113812 201006 113824
rect 317414 113812 317420 113824
rect 201000 113784 317420 113812
rect 201000 113772 201006 113784
rect 317414 113772 317420 113784
rect 317472 113772 317478 113824
rect 79686 113636 79692 113688
rect 79744 113676 79750 113688
rect 86862 113676 86868 113688
rect 79744 113648 86868 113676
rect 79744 113636 79750 113648
rect 86862 113636 86868 113648
rect 86920 113636 86926 113688
rect 70302 113568 70308 113620
rect 70360 113608 70366 113620
rect 72326 113608 72332 113620
rect 70360 113580 72332 113608
rect 70360 113568 70366 113580
rect 72326 113568 72332 113580
rect 72384 113568 72390 113620
rect 72436 113580 77294 113608
rect 67542 113500 67548 113552
rect 67600 113540 67606 113552
rect 72436 113540 72464 113580
rect 67600 113512 72464 113540
rect 77266 113540 77294 113580
rect 169110 113540 169116 113552
rect 77266 113512 169116 113540
rect 67600 113500 67606 113512
rect 169110 113500 169116 113512
rect 169168 113500 169174 113552
rect 72326 113432 72332 113484
rect 72384 113472 72390 113484
rect 162302 113472 162308 113484
rect 72384 113444 162308 113472
rect 72384 113432 72390 113444
rect 162302 113432 162308 113444
rect 162360 113432 162366 113484
rect 69382 113364 69388 113416
rect 69440 113404 69446 113416
rect 164970 113404 164976 113416
rect 69440 113376 164976 113404
rect 69440 113364 69446 113376
rect 164970 113364 164976 113376
rect 165028 113364 165034 113416
rect 68554 113296 68560 113348
rect 68612 113336 68618 113348
rect 165522 113336 165528 113348
rect 68612 113308 165528 113336
rect 68612 113296 68618 113308
rect 165522 113296 165528 113308
rect 165580 113296 165586 113348
rect 64506 113228 64512 113280
rect 64564 113268 64570 113280
rect 165338 113268 165344 113280
rect 64564 113240 165344 113268
rect 64564 113228 64570 113240
rect 165338 113228 165344 113240
rect 165396 113228 165402 113280
rect 200298 113268 200304 113280
rect 200132 113240 200304 113268
rect 166902 113160 166908 113212
rect 166960 113200 166966 113212
rect 169294 113200 169300 113212
rect 166960 113172 169300 113200
rect 166960 113160 166966 113172
rect 169294 113160 169300 113172
rect 169352 113160 169358 113212
rect 200132 112872 200160 113240
rect 200298 113228 200304 113240
rect 200356 113228 200362 113280
rect 200206 113160 200212 113212
rect 200264 113160 200270 113212
rect 200224 112872 200252 113160
rect 202230 113092 202236 113144
rect 202288 113132 202294 113144
rect 229922 113132 229928 113144
rect 202288 113104 229928 113132
rect 202288 113092 202294 113104
rect 229922 113092 229928 113104
rect 229980 113092 229986 113144
rect 200114 112820 200120 112872
rect 200172 112820 200178 112872
rect 200206 112820 200212 112872
rect 200264 112820 200270 112872
rect 69474 112480 69480 112532
rect 69532 112520 69538 112532
rect 137922 112520 137928 112532
rect 69532 112492 137928 112520
rect 69532 112480 69538 112492
rect 137922 112480 137928 112492
rect 137980 112480 137986 112532
rect 71590 112412 71596 112464
rect 71648 112452 71654 112464
rect 166902 112452 166908 112464
rect 71648 112424 166908 112452
rect 71648 112412 71654 112424
rect 166902 112412 166908 112424
rect 166960 112412 166966 112464
rect 67910 112344 67916 112396
rect 67968 112384 67974 112396
rect 157978 112384 157984 112396
rect 67968 112356 157984 112384
rect 67968 112344 67974 112356
rect 157978 112344 157984 112356
rect 158036 112344 158042 112396
rect 68738 112276 68744 112328
rect 68796 112316 68802 112328
rect 158714 112316 158720 112328
rect 68796 112288 158720 112316
rect 68796 112276 68802 112288
rect 158714 112276 158720 112288
rect 158772 112276 158778 112328
rect 69658 112208 69664 112260
rect 69716 112248 69722 112260
rect 162210 112248 162216 112260
rect 69716 112220 162216 112248
rect 69716 112208 69722 112220
rect 162210 112208 162216 112220
rect 162268 112208 162274 112260
rect 68462 112140 68468 112192
rect 68520 112180 68526 112192
rect 162118 112180 162124 112192
rect 68520 112152 162124 112180
rect 68520 112140 68526 112152
rect 162118 112140 162124 112152
rect 162176 112140 162182 112192
rect 67082 112072 67088 112124
rect 67140 112112 67146 112124
rect 162762 112112 162768 112124
rect 67140 112084 162768 112112
rect 67140 112072 67146 112084
rect 162762 112072 162768 112084
rect 162820 112072 162826 112124
rect 65518 112004 65524 112056
rect 65576 112044 65582 112056
rect 75178 112044 75184 112056
rect 65576 112016 75184 112044
rect 65576 112004 65582 112016
rect 75178 112004 75184 112016
rect 75236 112004 75242 112056
rect 75638 112004 75644 112056
rect 75696 112044 75702 112056
rect 166994 112044 167000 112056
rect 75696 112016 167000 112044
rect 75696 112004 75702 112016
rect 166994 112004 167000 112016
rect 167052 112004 167058 112056
rect 70026 111936 70032 111988
rect 70084 111976 70090 111988
rect 169386 111976 169392 111988
rect 70084 111948 75132 111976
rect 70084 111936 70090 111948
rect 67082 111868 67088 111920
rect 67140 111908 67146 111920
rect 67266 111908 67272 111920
rect 67140 111880 67272 111908
rect 67140 111868 67146 111880
rect 67266 111868 67272 111880
rect 67324 111868 67330 111920
rect 67818 111868 67824 111920
rect 67876 111908 67882 111920
rect 68462 111908 68468 111920
rect 67876 111880 68468 111908
rect 67876 111868 67882 111880
rect 68462 111868 68468 111880
rect 68520 111868 68526 111920
rect 68922 111868 68928 111920
rect 68980 111908 68986 111920
rect 70670 111908 70676 111920
rect 68980 111880 70676 111908
rect 68980 111868 68986 111880
rect 70670 111868 70676 111880
rect 70728 111908 70734 111920
rect 71590 111908 71596 111920
rect 70728 111880 71596 111908
rect 70728 111868 70734 111880
rect 71590 111868 71596 111880
rect 71648 111868 71654 111920
rect 75104 111908 75132 111948
rect 75380 111948 169392 111976
rect 75380 111908 75408 111948
rect 169386 111936 169392 111948
rect 169444 111936 169450 111988
rect 75104 111880 75408 111908
rect 75454 111868 75460 111920
rect 75512 111908 75518 111920
rect 101582 111908 101588 111920
rect 75512 111880 101588 111908
rect 75512 111868 75518 111880
rect 101582 111868 101588 111880
rect 101640 111868 101646 111920
rect 3418 111800 3424 111852
rect 3476 111840 3482 111852
rect 100754 111840 100760 111852
rect 3476 111812 100760 111840
rect 3476 111800 3482 111812
rect 100754 111800 100760 111812
rect 100812 111800 100818 111852
rect 158714 111800 158720 111852
rect 158772 111840 158778 111852
rect 159358 111840 159364 111852
rect 158772 111812 159364 111840
rect 158772 111800 158778 111812
rect 159358 111800 159364 111812
rect 159416 111800 159422 111852
rect 169386 111800 169392 111852
rect 169444 111840 169450 111852
rect 169662 111840 169668 111852
rect 169444 111812 169668 111840
rect 169444 111800 169450 111812
rect 169662 111800 169668 111812
rect 169720 111800 169726 111852
rect 63402 111732 63408 111784
rect 63460 111772 63466 111784
rect 68922 111772 68928 111784
rect 63460 111744 68928 111772
rect 63460 111732 63466 111744
rect 68922 111732 68928 111744
rect 68980 111732 68986 111784
rect 69290 111732 69296 111784
rect 69348 111772 69354 111784
rect 70302 111772 70308 111784
rect 69348 111744 70308 111772
rect 69348 111732 69354 111744
rect 70302 111732 70308 111744
rect 70360 111732 70366 111784
rect 108942 111732 108948 111784
rect 109000 111772 109006 111784
rect 111518 111772 111524 111784
rect 109000 111744 111524 111772
rect 109000 111732 109006 111744
rect 111518 111732 111524 111744
rect 111576 111772 111582 111784
rect 165246 111772 165252 111784
rect 111576 111744 165252 111772
rect 111576 111732 111582 111744
rect 165246 111732 165252 111744
rect 165304 111732 165310 111784
rect 69198 111664 69204 111716
rect 69256 111704 69262 111716
rect 69842 111704 69848 111716
rect 69256 111676 69848 111704
rect 69256 111664 69262 111676
rect 69842 111664 69848 111676
rect 69900 111704 69906 111716
rect 75638 111704 75644 111716
rect 69900 111676 75644 111704
rect 69900 111664 69906 111676
rect 75638 111664 75644 111676
rect 75696 111664 75702 111716
rect 105722 111664 105728 111716
rect 105780 111704 105786 111716
rect 119982 111704 119988 111716
rect 105780 111676 119988 111704
rect 105780 111664 105786 111676
rect 119982 111664 119988 111676
rect 120040 111704 120046 111716
rect 166442 111704 166448 111716
rect 120040 111676 166448 111704
rect 120040 111664 120046 111676
rect 166442 111664 166448 111676
rect 166500 111664 166506 111716
rect 108206 110508 108212 110560
rect 108264 110548 108270 110560
rect 108574 110548 108580 110560
rect 108264 110520 108580 110548
rect 108264 110508 108270 110520
rect 108574 110508 108580 110520
rect 108632 110508 108638 110560
rect 70302 110440 70308 110492
rect 70360 110480 70366 110492
rect 169478 110480 169484 110492
rect 70360 110452 169484 110480
rect 70360 110440 70366 110452
rect 169478 110440 169484 110452
rect 169536 110440 169542 110492
rect 108942 110372 108948 110424
rect 109000 110412 109006 110424
rect 165154 110412 165160 110424
rect 109000 110384 165160 110412
rect 109000 110372 109006 110384
rect 165154 110372 165160 110384
rect 165212 110372 165218 110424
rect 202782 110372 202788 110424
rect 202840 110412 202846 110424
rect 204714 110412 204720 110424
rect 202840 110384 204720 110412
rect 202840 110372 202846 110384
rect 204714 110372 204720 110384
rect 204772 110372 204778 110424
rect 108574 110304 108580 110356
rect 108632 110344 108638 110356
rect 121270 110344 121276 110356
rect 108632 110316 121276 110344
rect 108632 110304 108638 110316
rect 121270 110304 121276 110316
rect 121328 110304 121334 110356
rect 150434 110304 150440 110356
rect 150492 110344 150498 110356
rect 166994 110344 167000 110356
rect 150492 110316 167000 110344
rect 150492 110304 150498 110316
rect 166994 110304 167000 110316
rect 167052 110304 167058 110356
rect 201862 109760 201868 109812
rect 201920 109800 201926 109812
rect 203150 109800 203156 109812
rect 201920 109772 203156 109800
rect 201920 109760 201926 109772
rect 203150 109760 203156 109772
rect 203208 109800 203214 109812
rect 267826 109800 267832 109812
rect 203208 109772 267832 109800
rect 203208 109760 203214 109772
rect 267826 109760 267832 109772
rect 267884 109760 267890 109812
rect 204714 109692 204720 109744
rect 204772 109732 204778 109744
rect 299566 109732 299572 109744
rect 204772 109704 299572 109732
rect 204772 109692 204778 109704
rect 299566 109692 299572 109704
rect 299624 109692 299630 109744
rect 107654 108944 107660 108996
rect 107712 108984 107718 108996
rect 109770 108984 109776 108996
rect 107712 108956 109776 108984
rect 107712 108944 107718 108956
rect 109770 108944 109776 108956
rect 109828 108944 109834 108996
rect 116854 108984 116860 108996
rect 113146 108956 116860 108984
rect 108022 108876 108028 108928
rect 108080 108916 108086 108928
rect 113146 108916 113174 108956
rect 116854 108944 116860 108956
rect 116912 108944 116918 108996
rect 200298 108944 200304 108996
rect 200356 108984 200362 108996
rect 200482 108984 200488 108996
rect 200356 108956 200488 108984
rect 200356 108944 200362 108956
rect 200482 108944 200488 108956
rect 200540 108984 200546 108996
rect 230566 108984 230572 108996
rect 200540 108956 230572 108984
rect 200540 108944 200546 108956
rect 230566 108944 230572 108956
rect 230624 108984 230630 108996
rect 231762 108984 231768 108996
rect 230624 108956 231768 108984
rect 230624 108944 230630 108956
rect 231762 108944 231768 108956
rect 231820 108944 231826 108996
rect 108080 108888 113174 108916
rect 108080 108876 108086 108888
rect 167546 108332 167552 108384
rect 167604 108372 167610 108384
rect 167914 108372 167920 108384
rect 167604 108344 167920 108372
rect 167604 108332 167610 108344
rect 167914 108332 167920 108344
rect 167972 108332 167978 108384
rect 231762 108264 231768 108316
rect 231820 108304 231826 108316
rect 336734 108304 336740 108316
rect 231820 108276 336740 108304
rect 231820 108264 231826 108276
rect 336734 108264 336740 108276
rect 336792 108264 336798 108316
rect 165522 107584 165528 107636
rect 165580 107624 165586 107636
rect 166994 107624 167000 107636
rect 165580 107596 167000 107624
rect 165580 107584 165586 107596
rect 166994 107584 167000 107596
rect 167052 107584 167058 107636
rect 202782 107584 202788 107636
rect 202840 107624 202846 107636
rect 205726 107624 205732 107636
rect 202840 107596 205732 107624
rect 202840 107584 202846 107596
rect 205726 107584 205732 107596
rect 205784 107624 205790 107636
rect 230474 107624 230480 107636
rect 205784 107596 230480 107624
rect 205784 107584 205790 107596
rect 230474 107584 230480 107596
rect 230532 107624 230538 107636
rect 231762 107624 231768 107636
rect 230532 107596 231768 107624
rect 230532 107584 230538 107596
rect 231762 107584 231768 107596
rect 231820 107584 231826 107636
rect 108942 107448 108948 107500
rect 109000 107488 109006 107500
rect 164786 107488 164792 107500
rect 109000 107460 164792 107488
rect 109000 107448 109006 107460
rect 164786 107448 164792 107460
rect 164844 107448 164850 107500
rect 231762 106904 231768 106956
rect 231820 106944 231826 106956
rect 347774 106944 347780 106956
rect 231820 106916 347780 106944
rect 231820 106904 231826 106916
rect 347774 106904 347780 106916
rect 347832 106904 347838 106956
rect 108942 106632 108948 106684
rect 109000 106672 109006 106684
rect 112990 106672 112996 106684
rect 109000 106644 112996 106672
rect 109000 106632 109006 106644
rect 112990 106632 112996 106644
rect 113048 106632 113054 106684
rect 132494 106292 132500 106344
rect 132552 106332 132558 106344
rect 166994 106332 167000 106344
rect 132552 106304 167000 106332
rect 132552 106292 132558 106304
rect 166994 106292 167000 106304
rect 167052 106292 167058 106344
rect 108942 106224 108948 106276
rect 109000 106264 109006 106276
rect 165062 106264 165068 106276
rect 109000 106236 165068 106264
rect 109000 106224 109006 106236
rect 165062 106224 165068 106236
rect 165120 106224 165126 106276
rect 165338 106224 165344 106276
rect 165396 106264 165402 106276
rect 167914 106264 167920 106276
rect 165396 106236 167920 106264
rect 165396 106224 165402 106236
rect 167914 106224 167920 106236
rect 167972 106224 167978 106276
rect 201862 105544 201868 105596
rect 201920 105584 201926 105596
rect 230658 105584 230664 105596
rect 201920 105556 230664 105584
rect 201920 105544 201926 105556
rect 230658 105544 230664 105556
rect 230716 105544 230722 105596
rect 64506 104796 64512 104848
rect 64564 104836 64570 104848
rect 67634 104836 67640 104848
rect 64564 104808 67640 104836
rect 64564 104796 64570 104808
rect 67634 104796 67640 104808
rect 67692 104796 67698 104848
rect 108022 104796 108028 104848
rect 108080 104836 108086 104848
rect 119890 104836 119896 104848
rect 108080 104808 119896 104836
rect 108080 104796 108086 104808
rect 119890 104796 119896 104808
rect 119948 104796 119954 104848
rect 167454 104796 167460 104848
rect 167512 104836 167518 104848
rect 169202 104836 169208 104848
rect 167512 104808 169208 104836
rect 167512 104796 167518 104808
rect 169202 104796 169208 104808
rect 169260 104796 169266 104848
rect 200758 104116 200764 104168
rect 200816 104156 200822 104168
rect 289814 104156 289820 104168
rect 200816 104128 289820 104156
rect 200816 104116 200822 104128
rect 289814 104116 289820 104128
rect 289872 104116 289878 104168
rect 64782 103436 64788 103488
rect 64840 103476 64846 103488
rect 67634 103476 67640 103488
rect 64840 103448 67640 103476
rect 64840 103436 64846 103448
rect 67634 103436 67640 103448
rect 67692 103436 67698 103488
rect 108942 103436 108948 103488
rect 109000 103476 109006 103488
rect 147030 103476 147036 103488
rect 109000 103448 147036 103476
rect 109000 103436 109006 103448
rect 147030 103436 147036 103448
rect 147088 103436 147094 103488
rect 162026 103436 162032 103488
rect 162084 103476 162090 103488
rect 166994 103476 167000 103488
rect 162084 103448 167000 103476
rect 162084 103436 162090 103448
rect 166994 103436 167000 103448
rect 167052 103436 167058 103488
rect 108206 103368 108212 103420
rect 108264 103408 108270 103420
rect 121362 103408 121368 103420
rect 108264 103380 121368 103408
rect 108264 103368 108270 103380
rect 121362 103368 121368 103380
rect 121420 103368 121426 103420
rect 203702 102756 203708 102808
rect 203760 102796 203766 102808
rect 255314 102796 255320 102808
rect 203760 102768 255320 102796
rect 203760 102756 203766 102768
rect 255314 102756 255320 102768
rect 255372 102756 255378 102808
rect 162762 102076 162768 102128
rect 162820 102116 162826 102128
rect 166994 102116 167000 102128
rect 162820 102088 167000 102116
rect 162820 102076 162826 102088
rect 166994 102076 167000 102088
rect 167052 102076 167058 102128
rect 108942 102008 108948 102060
rect 109000 102048 109006 102060
rect 115290 102048 115296 102060
rect 109000 102020 115296 102048
rect 109000 102008 109006 102020
rect 115290 102008 115296 102020
rect 115348 102008 115354 102060
rect 108574 101736 108580 101788
rect 108632 101776 108638 101788
rect 108758 101776 108764 101788
rect 108632 101748 108764 101776
rect 108632 101736 108638 101748
rect 108758 101736 108764 101748
rect 108816 101736 108822 101788
rect 108758 101600 108764 101652
rect 108816 101640 108822 101652
rect 115382 101640 115388 101652
rect 108816 101612 115388 101640
rect 108816 101600 108822 101612
rect 115382 101600 115388 101612
rect 115440 101600 115446 101652
rect 66070 100648 66076 100700
rect 66128 100688 66134 100700
rect 67634 100688 67640 100700
rect 66128 100660 67640 100688
rect 66128 100648 66134 100660
rect 67634 100648 67640 100660
rect 67692 100648 67698 100700
rect 108942 100648 108948 100700
rect 109000 100688 109006 100700
rect 162578 100688 162584 100700
rect 109000 100660 162584 100688
rect 109000 100648 109006 100660
rect 162578 100648 162584 100660
rect 162636 100648 162642 100700
rect 163498 100648 163504 100700
rect 163556 100688 163562 100700
rect 167454 100688 167460 100700
rect 163556 100660 167460 100688
rect 163556 100648 163562 100660
rect 167454 100648 167460 100660
rect 167512 100648 167518 100700
rect 66162 100580 66168 100632
rect 66220 100620 66226 100632
rect 68278 100620 68284 100632
rect 66220 100592 68284 100620
rect 66220 100580 66226 100592
rect 68278 100580 68284 100592
rect 68336 100580 68342 100632
rect 108758 100580 108764 100632
rect 108816 100620 108822 100632
rect 159542 100620 159548 100632
rect 108816 100592 159548 100620
rect 108816 100580 108822 100592
rect 159542 100580 159548 100592
rect 159600 100580 159606 100632
rect 155218 100512 155224 100564
rect 155276 100552 155282 100564
rect 167086 100552 167092 100564
rect 155276 100524 167092 100552
rect 155276 100512 155282 100524
rect 167086 100512 167092 100524
rect 167144 100512 167150 100564
rect 202782 100036 202788 100088
rect 202840 100076 202846 100088
rect 208394 100076 208400 100088
rect 202840 100048 208400 100076
rect 202840 100036 202846 100048
rect 208394 100036 208400 100048
rect 208452 100076 208458 100088
rect 256694 100076 256700 100088
rect 208452 100048 256700 100076
rect 208452 100036 208458 100048
rect 256694 100036 256700 100048
rect 256752 100036 256758 100088
rect 201586 99968 201592 100020
rect 201644 100008 201650 100020
rect 204622 100008 204628 100020
rect 201644 99980 204628 100008
rect 201644 99968 201650 99980
rect 204622 99968 204628 99980
rect 204680 100008 204686 100020
rect 307846 100008 307852 100020
rect 204680 99980 307852 100008
rect 204680 99968 204686 99980
rect 307846 99968 307852 99980
rect 307904 99968 307910 100020
rect 258718 99356 258724 99408
rect 258776 99396 258782 99408
rect 580166 99396 580172 99408
rect 258776 99368 580172 99396
rect 258776 99356 258782 99368
rect 580166 99356 580172 99368
rect 580224 99356 580230 99408
rect 64322 99288 64328 99340
rect 64380 99328 64386 99340
rect 67634 99328 67640 99340
rect 64380 99300 67640 99328
rect 64380 99288 64386 99300
rect 67634 99288 67640 99300
rect 67692 99288 67698 99340
rect 107654 99288 107660 99340
rect 107712 99328 107718 99340
rect 162486 99328 162492 99340
rect 107712 99300 162492 99328
rect 107712 99288 107718 99300
rect 162486 99288 162492 99300
rect 162544 99288 162550 99340
rect 201586 99288 201592 99340
rect 201644 99328 201650 99340
rect 219434 99328 219440 99340
rect 201644 99300 219440 99328
rect 201644 99288 201650 99300
rect 219434 99288 219440 99300
rect 219492 99288 219498 99340
rect 107746 98608 107752 98660
rect 107804 98648 107810 98660
rect 119614 98648 119620 98660
rect 107804 98620 119620 98648
rect 107804 98608 107810 98620
rect 119614 98608 119620 98620
rect 119672 98608 119678 98660
rect 65978 97928 65984 97980
rect 66036 97968 66042 97980
rect 67634 97968 67640 97980
rect 66036 97940 67640 97968
rect 66036 97928 66042 97940
rect 67634 97928 67640 97940
rect 67692 97928 67698 97980
rect 107654 97928 107660 97980
rect 107712 97968 107718 97980
rect 121086 97968 121092 97980
rect 107712 97940 121092 97968
rect 107712 97928 107718 97940
rect 121086 97928 121092 97940
rect 121144 97928 121150 97980
rect 165522 97928 165528 97980
rect 165580 97968 165586 97980
rect 166350 97968 166356 97980
rect 165580 97940 166356 97968
rect 165580 97928 165586 97940
rect 166350 97928 166356 97940
rect 166408 97928 166414 97980
rect 162210 97860 162216 97912
rect 162268 97900 162274 97912
rect 167178 97900 167184 97912
rect 162268 97872 167184 97900
rect 162268 97860 162274 97872
rect 167178 97860 167184 97872
rect 167236 97860 167242 97912
rect 108390 96636 108396 96688
rect 108448 96676 108454 96688
rect 165522 96676 165528 96688
rect 108448 96648 165528 96676
rect 108448 96636 108454 96648
rect 165522 96636 165528 96648
rect 165580 96636 165586 96688
rect 64230 96568 64236 96620
rect 64288 96608 64294 96620
rect 67634 96608 67640 96620
rect 64288 96580 67640 96608
rect 64288 96568 64294 96580
rect 67634 96568 67640 96580
rect 67692 96568 67698 96620
rect 107838 96568 107844 96620
rect 107896 96608 107902 96620
rect 119706 96608 119712 96620
rect 107896 96580 119712 96608
rect 107896 96568 107902 96580
rect 119706 96568 119712 96580
rect 119764 96568 119770 96620
rect 159358 96568 159364 96620
rect 159416 96608 159422 96620
rect 168834 96608 168840 96620
rect 159416 96580 168840 96608
rect 159416 96568 159422 96580
rect 168834 96568 168840 96580
rect 168892 96568 168898 96620
rect 66622 96500 66628 96552
rect 66680 96540 66686 96552
rect 69198 96540 69204 96552
rect 66680 96512 69204 96540
rect 66680 96500 66686 96512
rect 69198 96500 69204 96512
rect 69256 96500 69262 96552
rect 107654 96500 107660 96552
rect 107712 96540 107718 96552
rect 119246 96540 119252 96552
rect 107712 96512 119252 96540
rect 107712 96500 107718 96512
rect 119246 96500 119252 96512
rect 119304 96500 119310 96552
rect 202138 95888 202144 95940
rect 202196 95928 202202 95940
rect 203058 95928 203064 95940
rect 202196 95900 203064 95928
rect 202196 95888 202202 95900
rect 203058 95888 203064 95900
rect 203116 95928 203122 95940
rect 260834 95928 260840 95940
rect 203116 95900 260840 95928
rect 203116 95888 203122 95900
rect 260834 95888 260840 95900
rect 260892 95888 260898 95940
rect 107746 95208 107752 95260
rect 107804 95248 107810 95260
rect 166442 95248 166448 95260
rect 107804 95220 166448 95248
rect 107804 95208 107810 95220
rect 166442 95208 166448 95220
rect 166500 95208 166506 95260
rect 201402 95208 201408 95260
rect 201460 95248 201466 95260
rect 324314 95248 324320 95260
rect 201460 95220 324320 95248
rect 201460 95208 201466 95220
rect 324314 95208 324320 95220
rect 324372 95208 324378 95260
rect 107654 95140 107660 95192
rect 107712 95180 107718 95192
rect 120074 95180 120080 95192
rect 107712 95152 120080 95180
rect 107712 95140 107718 95152
rect 120074 95140 120080 95152
rect 120132 95180 120138 95192
rect 120626 95180 120632 95192
rect 120132 95152 120632 95180
rect 120132 95140 120138 95152
rect 120626 95140 120632 95152
rect 120684 95140 120690 95192
rect 137922 95140 137928 95192
rect 137980 95180 137986 95192
rect 166994 95180 167000 95192
rect 137980 95152 167000 95180
rect 137980 95140 137986 95152
rect 166994 95140 167000 95152
rect 167052 95140 167058 95192
rect 120074 94528 120080 94580
rect 120132 94568 120138 94580
rect 166350 94568 166356 94580
rect 120132 94540 166356 94568
rect 120132 94528 120138 94540
rect 166350 94528 166356 94540
rect 166408 94528 166414 94580
rect 107654 94460 107660 94512
rect 107712 94500 107718 94512
rect 119982 94500 119988 94512
rect 107712 94472 119988 94500
rect 107712 94460 107718 94472
rect 119982 94460 119988 94472
rect 120040 94500 120046 94512
rect 166534 94500 166540 94512
rect 120040 94472 166540 94500
rect 120040 94460 120046 94472
rect 166534 94460 166540 94472
rect 166592 94460 166598 94512
rect 202782 94460 202788 94512
rect 202840 94500 202846 94512
rect 204530 94500 204536 94512
rect 202840 94472 204536 94500
rect 202840 94460 202846 94472
rect 204530 94460 204536 94472
rect 204588 94500 204594 94512
rect 296714 94500 296720 94512
rect 204588 94472 296720 94500
rect 204588 94460 204594 94472
rect 296714 94460 296720 94472
rect 296772 94460 296778 94512
rect 64690 93780 64696 93832
rect 64748 93820 64754 93832
rect 67634 93820 67640 93832
rect 64748 93792 67640 93820
rect 64748 93780 64754 93792
rect 67634 93780 67640 93792
rect 67692 93780 67698 93832
rect 107746 93780 107752 93832
rect 107804 93820 107810 93832
rect 162394 93820 162400 93832
rect 107804 93792 162400 93820
rect 107804 93780 107810 93792
rect 162394 93780 162400 93792
rect 162452 93780 162458 93832
rect 107654 93712 107660 93764
rect 107712 93752 107718 93764
rect 120902 93752 120908 93764
rect 107712 93724 120908 93752
rect 107712 93712 107718 93724
rect 120902 93712 120908 93724
rect 120960 93712 120966 93764
rect 64414 92420 64420 92472
rect 64472 92460 64478 92472
rect 67634 92460 67640 92472
rect 64472 92432 67640 92460
rect 64472 92420 64478 92432
rect 67634 92420 67640 92432
rect 67692 92420 67698 92472
rect 65702 92352 65708 92404
rect 65760 92392 65766 92404
rect 68094 92392 68100 92404
rect 65760 92364 68100 92392
rect 65760 92352 65766 92364
rect 68094 92352 68100 92364
rect 68152 92352 68158 92404
rect 107746 91740 107752 91792
rect 107804 91780 107810 91792
rect 122282 91780 122288 91792
rect 107804 91752 122288 91780
rect 107804 91740 107810 91752
rect 122282 91740 122288 91752
rect 122340 91740 122346 91792
rect 164970 90992 164976 91044
rect 165028 91032 165034 91044
rect 167638 91032 167644 91044
rect 165028 91004 167644 91032
rect 165028 90992 165034 91004
rect 167638 90992 167644 91004
rect 167696 90992 167702 91044
rect 201770 90788 201776 90840
rect 201828 90828 201834 90840
rect 204438 90828 204444 90840
rect 201828 90800 204444 90828
rect 201828 90788 201834 90800
rect 204438 90788 204444 90800
rect 204496 90788 204502 90840
rect 108022 90380 108028 90432
rect 108080 90420 108086 90432
rect 120810 90420 120816 90432
rect 108080 90392 120816 90420
rect 108080 90380 108086 90392
rect 120810 90380 120816 90392
rect 120868 90380 120874 90432
rect 107654 90312 107660 90364
rect 107712 90352 107718 90364
rect 119338 90352 119344 90364
rect 107712 90324 119344 90352
rect 107712 90312 107718 90324
rect 119338 90312 119344 90324
rect 119396 90352 119402 90364
rect 165062 90352 165068 90364
rect 119396 90324 165068 90352
rect 119396 90312 119402 90324
rect 165062 90312 165068 90324
rect 165120 90312 165126 90364
rect 204438 90312 204444 90364
rect 204496 90352 204502 90364
rect 346394 90352 346400 90364
rect 204496 90324 346400 90352
rect 204496 90312 204502 90324
rect 346394 90312 346400 90324
rect 346452 90312 346458 90364
rect 201770 90040 201776 90092
rect 201828 90080 201834 90092
rect 208394 90080 208400 90092
rect 201828 90052 208400 90080
rect 201828 90040 201834 90052
rect 208394 90040 208400 90052
rect 208452 90040 208458 90092
rect 107102 89700 107108 89752
rect 107160 89740 107166 89752
rect 166994 89740 167000 89752
rect 107160 89712 167000 89740
rect 107160 89700 107166 89712
rect 166994 89700 167000 89712
rect 167052 89700 167058 89752
rect 157978 89632 157984 89684
rect 158036 89672 158042 89684
rect 167178 89672 167184 89684
rect 158036 89644 167184 89672
rect 158036 89632 158042 89644
rect 167178 89632 167184 89644
rect 167236 89632 167242 89684
rect 202506 89632 202512 89684
rect 202564 89672 202570 89684
rect 229094 89672 229100 89684
rect 202564 89644 229100 89672
rect 202564 89632 202570 89644
rect 229094 89632 229100 89644
rect 229152 89672 229158 89684
rect 230382 89672 230388 89684
rect 229152 89644 230388 89672
rect 229152 89632 229158 89644
rect 230382 89632 230388 89644
rect 230440 89632 230446 89684
rect 108574 88952 108580 89004
rect 108632 88992 108638 89004
rect 166626 88992 166632 89004
rect 108632 88964 166632 88992
rect 108632 88952 108638 88964
rect 166626 88952 166632 88964
rect 166684 88952 166690 89004
rect 230382 88952 230388 89004
rect 230440 88992 230446 89004
rect 329834 88992 329840 89004
rect 230440 88964 329840 88992
rect 230440 88952 230446 88964
rect 329834 88952 329840 88964
rect 329892 88952 329898 89004
rect 66898 88476 66904 88528
rect 66956 88516 66962 88528
rect 68462 88516 68468 88528
rect 66956 88488 68468 88516
rect 66956 88476 66962 88488
rect 68462 88476 68468 88488
rect 68520 88476 68526 88528
rect 107286 88340 107292 88392
rect 107344 88380 107350 88392
rect 166994 88380 167000 88392
rect 107344 88352 167000 88380
rect 107344 88340 107350 88352
rect 166994 88340 167000 88352
rect 167052 88340 167058 88392
rect 108942 88272 108948 88324
rect 109000 88312 109006 88324
rect 119522 88312 119528 88324
rect 109000 88284 119528 88312
rect 109000 88272 109006 88284
rect 119522 88272 119528 88284
rect 119580 88272 119586 88324
rect 162302 88272 162308 88324
rect 162360 88312 162366 88324
rect 167086 88312 167092 88324
rect 162360 88284 167092 88312
rect 162360 88272 162366 88284
rect 167086 88272 167092 88284
rect 167144 88272 167150 88324
rect 202506 88272 202512 88324
rect 202564 88312 202570 88324
rect 226334 88312 226340 88324
rect 202564 88284 226340 88312
rect 202564 88272 202570 88284
rect 226334 88272 226340 88284
rect 226392 88312 226398 88324
rect 226794 88312 226800 88324
rect 226392 88284 226800 88312
rect 226392 88272 226398 88284
rect 226794 88272 226800 88284
rect 226852 88272 226858 88324
rect 226794 87592 226800 87644
rect 226852 87632 226858 87644
rect 316034 87632 316040 87644
rect 226852 87604 316040 87632
rect 226852 87592 226858 87604
rect 316034 87592 316040 87604
rect 316092 87592 316098 87644
rect 3418 86980 3424 87032
rect 3476 87020 3482 87032
rect 68094 87020 68100 87032
rect 3476 86992 68100 87020
rect 3476 86980 3482 86992
rect 68094 86980 68100 86992
rect 68152 86980 68158 87032
rect 67450 86912 67456 86964
rect 67508 86952 67514 86964
rect 67910 86952 67916 86964
rect 67508 86924 67916 86952
rect 67508 86912 67514 86924
rect 67910 86912 67916 86924
rect 67968 86912 67974 86964
rect 108942 86912 108948 86964
rect 109000 86952 109006 86964
rect 119430 86952 119436 86964
rect 109000 86924 119436 86952
rect 109000 86912 109006 86924
rect 119430 86912 119436 86924
rect 119488 86912 119494 86964
rect 164142 86912 164148 86964
rect 164200 86952 164206 86964
rect 164878 86952 164884 86964
rect 164200 86924 164884 86952
rect 164200 86912 164206 86924
rect 164878 86912 164884 86924
rect 164936 86912 164942 86964
rect 202506 86912 202512 86964
rect 202564 86952 202570 86964
rect 227806 86952 227812 86964
rect 202564 86924 227812 86952
rect 202564 86912 202570 86924
rect 227806 86912 227812 86924
rect 227864 86912 227870 86964
rect 227806 86232 227812 86284
rect 227864 86272 227870 86284
rect 238754 86272 238760 86284
rect 227864 86244 238760 86272
rect 227864 86232 227870 86244
rect 238754 86232 238760 86244
rect 238812 86232 238818 86284
rect 200114 86096 200120 86148
rect 200172 86096 200178 86148
rect 111058 85620 111064 85672
rect 111116 85660 111122 85672
rect 164142 85660 164148 85672
rect 111116 85632 164148 85660
rect 111116 85620 111122 85632
rect 164142 85620 164148 85632
rect 164200 85620 164206 85672
rect 107194 85552 107200 85604
rect 107252 85592 107258 85604
rect 166994 85592 167000 85604
rect 107252 85564 167000 85592
rect 107252 85552 107258 85564
rect 166994 85552 167000 85564
rect 167052 85552 167058 85604
rect 200132 85536 200160 86096
rect 233878 85552 233884 85604
rect 233936 85592 233942 85604
rect 580166 85592 580172 85604
rect 233936 85564 580172 85592
rect 233936 85552 233942 85564
rect 580166 85552 580172 85564
rect 580224 85552 580230 85604
rect 108206 85484 108212 85536
rect 108264 85524 108270 85536
rect 144822 85524 144828 85536
rect 108264 85496 144828 85524
rect 108264 85484 108270 85496
rect 144822 85484 144828 85496
rect 144880 85484 144886 85536
rect 162118 85484 162124 85536
rect 162176 85524 162182 85536
rect 167086 85524 167092 85536
rect 162176 85496 167092 85524
rect 162176 85484 162182 85496
rect 167086 85484 167092 85496
rect 167144 85484 167150 85536
rect 200114 85484 200120 85536
rect 200172 85484 200178 85536
rect 3326 84804 3332 84856
rect 3384 84844 3390 84856
rect 67634 84844 67640 84856
rect 3384 84816 67640 84844
rect 3384 84804 3390 84816
rect 67634 84804 67640 84816
rect 67692 84844 67698 84856
rect 67818 84844 67824 84856
rect 67692 84816 67824 84844
rect 67692 84804 67698 84816
rect 67818 84804 67824 84816
rect 67876 84804 67882 84856
rect 109218 84804 109224 84856
rect 109276 84844 109282 84856
rect 122190 84844 122196 84856
rect 109276 84816 122196 84844
rect 109276 84804 109282 84816
rect 122190 84804 122196 84816
rect 122248 84804 122254 84856
rect 144822 84804 144828 84856
rect 144880 84844 144886 84856
rect 164878 84844 164884 84856
rect 144880 84816 164884 84844
rect 144880 84804 144886 84816
rect 164878 84804 164884 84816
rect 164936 84804 164942 84856
rect 202690 84804 202696 84856
rect 202748 84844 202754 84856
rect 203242 84844 203248 84856
rect 202748 84816 203248 84844
rect 202748 84804 202754 84816
rect 203242 84804 203248 84816
rect 203300 84844 203306 84856
rect 215202 84844 215208 84856
rect 203300 84816 215208 84844
rect 203300 84804 203306 84816
rect 215202 84804 215208 84816
rect 215260 84844 215266 84856
rect 277394 84844 277400 84856
rect 215260 84816 277400 84844
rect 215260 84804 215266 84816
rect 277394 84804 277400 84816
rect 277452 84804 277458 84856
rect 202690 84192 202696 84244
rect 202748 84232 202754 84244
rect 203058 84232 203064 84244
rect 202748 84204 203064 84232
rect 202748 84192 202754 84204
rect 203058 84192 203064 84204
rect 203116 84232 203122 84244
rect 332594 84232 332600 84244
rect 203116 84204 332600 84232
rect 203116 84192 203122 84204
rect 332594 84192 332600 84204
rect 332652 84192 332658 84244
rect 108942 84124 108948 84176
rect 109000 84164 109006 84176
rect 157242 84164 157248 84176
rect 109000 84136 157248 84164
rect 109000 84124 109006 84136
rect 157242 84124 157248 84136
rect 157300 84124 157306 84176
rect 157242 83512 157248 83564
rect 157300 83552 157306 83564
rect 166810 83552 166816 83564
rect 157300 83524 166816 83552
rect 157300 83512 157306 83524
rect 166810 83512 166816 83524
rect 166868 83512 166874 83564
rect 155862 83444 155868 83496
rect 155920 83484 155926 83496
rect 166994 83484 167000 83496
rect 155920 83456 167000 83484
rect 155920 83444 155926 83456
rect 166994 83444 167000 83456
rect 167052 83444 167058 83496
rect 203150 83444 203156 83496
rect 203208 83484 203214 83496
rect 224862 83484 224868 83496
rect 203208 83456 224868 83484
rect 203208 83444 203214 83456
rect 224862 83444 224868 83456
rect 224920 83484 224926 83496
rect 331214 83484 331220 83496
rect 224920 83456 331220 83484
rect 224920 83444 224926 83456
rect 331214 83444 331220 83456
rect 331272 83444 331278 83496
rect 117222 82832 117228 82884
rect 117280 82872 117286 82884
rect 162118 82872 162124 82884
rect 117280 82844 162124 82872
rect 117280 82832 117286 82844
rect 162118 82832 162124 82844
rect 162176 82832 162182 82884
rect 108942 82764 108948 82816
rect 109000 82804 109006 82816
rect 117240 82804 117268 82832
rect 109000 82776 117268 82804
rect 109000 82764 109006 82776
rect 67358 82356 67364 82408
rect 67416 82396 67422 82408
rect 68462 82396 68468 82408
rect 67416 82368 68468 82396
rect 67416 82356 67422 82368
rect 68462 82356 68468 82368
rect 68520 82356 68526 82408
rect 108850 82084 108856 82136
rect 108908 82124 108914 82136
rect 166902 82124 166908 82136
rect 108908 82096 166908 82124
rect 108908 82084 108914 82096
rect 166902 82084 166908 82096
rect 166960 82084 166966 82136
rect 107378 81404 107384 81456
rect 107436 81444 107442 81456
rect 166994 81444 167000 81456
rect 107436 81416 167000 81444
rect 107436 81404 107442 81416
rect 166994 81404 167000 81416
rect 167052 81404 167058 81456
rect 108942 81336 108948 81388
rect 109000 81376 109006 81388
rect 116762 81376 116768 81388
rect 109000 81348 116768 81376
rect 109000 81336 109006 81348
rect 116762 81336 116768 81348
rect 116820 81336 116826 81388
rect 108850 81268 108856 81320
rect 108908 81308 108914 81320
rect 112530 81308 112536 81320
rect 108908 81280 112536 81308
rect 108908 81268 108914 81280
rect 112530 81268 112536 81280
rect 112588 81268 112594 81320
rect 151722 80656 151728 80708
rect 151780 80696 151786 80708
rect 166994 80696 167000 80708
rect 151780 80668 167000 80696
rect 151780 80656 151786 80668
rect 166994 80656 167000 80668
rect 167052 80656 167058 80708
rect 107746 79976 107752 80028
rect 107804 80016 107810 80028
rect 120718 80016 120724 80028
rect 107804 79988 120724 80016
rect 107804 79976 107810 79988
rect 120718 79976 120724 79988
rect 120776 79976 120782 80028
rect 166166 79296 166172 79348
rect 166224 79336 166230 79348
rect 166718 79336 166724 79348
rect 166224 79308 166724 79336
rect 166224 79296 166230 79308
rect 166718 79296 166724 79308
rect 166776 79296 166782 79348
rect 202782 79296 202788 79348
rect 202840 79336 202846 79348
rect 203334 79336 203340 79348
rect 202840 79308 203340 79336
rect 202840 79296 202846 79308
rect 203334 79296 203340 79308
rect 203392 79336 203398 79348
rect 217962 79336 217968 79348
rect 203392 79308 217968 79336
rect 203392 79296 203398 79308
rect 217962 79296 217968 79308
rect 218020 79336 218026 79348
rect 241514 79336 241520 79348
rect 218020 79308 241520 79336
rect 218020 79296 218026 79308
rect 241514 79296 241520 79308
rect 241572 79296 241578 79348
rect 108666 79228 108672 79280
rect 108724 79268 108730 79280
rect 111886 79268 111892 79280
rect 108724 79240 111892 79268
rect 108724 79228 108730 79240
rect 111886 79228 111892 79240
rect 111944 79228 111950 79280
rect 118142 78752 118148 78804
rect 118200 78792 118206 78804
rect 118510 78792 118516 78804
rect 118200 78764 118516 78792
rect 118200 78752 118206 78764
rect 118510 78752 118516 78764
rect 118568 78792 118574 78804
rect 164970 78792 164976 78804
rect 118568 78764 164976 78792
rect 118568 78752 118574 78764
rect 164970 78752 164976 78764
rect 165028 78752 165034 78804
rect 165154 78752 165160 78804
rect 165212 78792 165218 78804
rect 166994 78792 167000 78804
rect 165212 78764 167000 78792
rect 165212 78752 165218 78764
rect 166994 78752 167000 78764
rect 167052 78752 167058 78804
rect 4798 78684 4804 78736
rect 4856 78724 4862 78736
rect 65978 78724 65984 78736
rect 4856 78696 65984 78724
rect 4856 78684 4862 78696
rect 65978 78684 65984 78696
rect 66036 78724 66042 78736
rect 67634 78724 67640 78736
rect 66036 78696 67640 78724
rect 66036 78684 66042 78696
rect 67634 78684 67640 78696
rect 67692 78684 67698 78736
rect 106918 78684 106924 78736
rect 106976 78724 106982 78736
rect 107930 78724 107936 78736
rect 106976 78696 107936 78724
rect 106976 78684 106982 78696
rect 107930 78684 107936 78696
rect 107988 78724 107994 78736
rect 166258 78724 166264 78736
rect 107988 78696 166264 78724
rect 107988 78684 107994 78696
rect 166258 78684 166264 78696
rect 166316 78684 166322 78736
rect 202782 78684 202788 78736
rect 202840 78724 202846 78736
rect 204438 78724 204444 78736
rect 202840 78696 204444 78724
rect 202840 78684 202846 78696
rect 204438 78684 204444 78696
rect 204496 78684 204502 78736
rect 65426 78616 65432 78668
rect 65484 78656 65490 78668
rect 66162 78656 66168 78668
rect 65484 78628 66168 78656
rect 65484 78616 65490 78628
rect 66162 78616 66168 78628
rect 66220 78616 66226 78668
rect 107746 78616 107752 78668
rect 107804 78656 107810 78668
rect 118142 78656 118148 78668
rect 107804 78628 118148 78656
rect 107804 78616 107810 78628
rect 118142 78616 118148 78628
rect 118200 78616 118206 78668
rect 65334 78548 65340 78600
rect 65392 78588 65398 78600
rect 66070 78588 66076 78600
rect 65392 78560 66076 78588
rect 65392 78548 65398 78560
rect 66070 78548 66076 78560
rect 66128 78588 66134 78600
rect 67634 78588 67640 78600
rect 66128 78560 67640 78588
rect 66128 78548 66134 78560
rect 67634 78548 67640 78560
rect 67692 78548 67698 78600
rect 66162 77596 66168 77648
rect 66220 77636 66226 77648
rect 67634 77636 67640 77648
rect 66220 77608 67640 77636
rect 66220 77596 66226 77608
rect 67634 77596 67640 77608
rect 67692 77596 67698 77648
rect 111610 77296 111616 77308
rect 110432 77268 111616 77296
rect 107746 77188 107752 77240
rect 107804 77228 107810 77240
rect 110432 77228 110460 77268
rect 111610 77256 111616 77268
rect 111668 77296 111674 77308
rect 162210 77296 162216 77308
rect 111668 77268 162216 77296
rect 111668 77256 111674 77268
rect 162210 77256 162216 77268
rect 162268 77256 162274 77308
rect 107804 77200 110460 77228
rect 107804 77188 107810 77200
rect 118142 76032 118148 76084
rect 118200 76072 118206 76084
rect 118602 76072 118608 76084
rect 118200 76044 118608 76072
rect 118200 76032 118206 76044
rect 118602 76032 118608 76044
rect 118660 76072 118666 76084
rect 162394 76072 162400 76084
rect 118660 76044 162400 76072
rect 118660 76032 118666 76044
rect 162394 76032 162400 76044
rect 162452 76032 162458 76084
rect 107838 75964 107844 76016
rect 107896 76004 107902 76016
rect 108114 76004 108120 76016
rect 107896 75976 108120 76004
rect 107896 75964 107902 75976
rect 108114 75964 108120 75976
rect 108172 76004 108178 76016
rect 162302 76004 162308 76016
rect 108172 75976 162308 76004
rect 108172 75964 108178 75976
rect 162302 75964 162308 75976
rect 162360 75964 162366 76016
rect 107746 75896 107752 75948
rect 107804 75936 107810 75948
rect 162854 75936 162860 75948
rect 107804 75908 162860 75936
rect 107804 75896 107810 75908
rect 162854 75896 162860 75908
rect 162912 75896 162918 75948
rect 201310 75896 201316 75948
rect 201368 75936 201374 75948
rect 253934 75936 253940 75948
rect 201368 75908 253940 75936
rect 201368 75896 201374 75908
rect 253934 75896 253940 75908
rect 253992 75896 253998 75948
rect 200942 75828 200948 75880
rect 201000 75868 201006 75880
rect 222838 75868 222844 75880
rect 201000 75840 222844 75868
rect 201000 75828 201006 75840
rect 222838 75828 222844 75840
rect 222896 75868 222902 75880
rect 223482 75868 223488 75880
rect 222896 75840 223488 75868
rect 222896 75828 222902 75840
rect 223482 75828 223488 75840
rect 223540 75828 223546 75880
rect 107838 75216 107844 75268
rect 107896 75256 107902 75268
rect 118142 75256 118148 75268
rect 107896 75228 118148 75256
rect 107896 75216 107902 75228
rect 118142 75216 118148 75228
rect 118200 75216 118206 75268
rect 107746 75148 107752 75200
rect 107804 75188 107810 75200
rect 111702 75188 111708 75200
rect 107804 75160 111708 75188
rect 107804 75148 107810 75160
rect 111702 75148 111708 75160
rect 111760 75188 111766 75200
rect 166718 75188 166724 75200
rect 111760 75160 166724 75188
rect 111760 75148 111766 75160
rect 166718 75148 166724 75160
rect 166776 75148 166782 75200
rect 223482 75148 223488 75200
rect 223540 75188 223546 75200
rect 302234 75188 302240 75200
rect 223540 75160 302240 75188
rect 223540 75148 223546 75160
rect 302234 75148 302240 75160
rect 302292 75148 302298 75200
rect 106182 74536 106188 74588
rect 106240 74576 106246 74588
rect 167086 74576 167092 74588
rect 106240 74548 167092 74576
rect 106240 74536 106246 74548
rect 167086 74536 167092 74548
rect 167144 74536 167150 74588
rect 200482 74536 200488 74588
rect 200540 74576 200546 74588
rect 339494 74576 339500 74588
rect 200540 74548 339500 74576
rect 200540 74536 200546 74548
rect 339494 74536 339500 74548
rect 339552 74536 339558 74588
rect 107746 74468 107752 74520
rect 107804 74508 107810 74520
rect 153102 74508 153108 74520
rect 107804 74480 153108 74508
rect 107804 74468 107810 74480
rect 153102 74468 153108 74480
rect 153160 74468 153166 74520
rect 201954 74468 201960 74520
rect 202012 74508 202018 74520
rect 221458 74508 221464 74520
rect 202012 74480 221464 74508
rect 202012 74468 202018 74480
rect 221458 74468 221464 74480
rect 221516 74468 221522 74520
rect 117958 73312 117964 73364
rect 118016 73352 118022 73364
rect 164786 73352 164792 73364
rect 118016 73324 164792 73352
rect 118016 73312 118022 73324
rect 164786 73312 164792 73324
rect 164844 73312 164850 73364
rect 165522 73244 165528 73296
rect 165580 73284 165586 73296
rect 167178 73284 167184 73296
rect 165580 73256 167184 73284
rect 165580 73244 165586 73256
rect 167178 73244 167184 73256
rect 167236 73244 167242 73296
rect 106090 73176 106096 73228
rect 106148 73216 106154 73228
rect 167086 73216 167092 73228
rect 106148 73188 167092 73216
rect 106148 73176 106154 73188
rect 167086 73176 167092 73188
rect 167144 73176 167150 73228
rect 107746 73108 107752 73160
rect 107804 73148 107810 73160
rect 117958 73148 117964 73160
rect 107804 73120 117964 73148
rect 107804 73108 107810 73120
rect 117958 73108 117964 73120
rect 118016 73108 118022 73160
rect 66714 72428 66720 72480
rect 66772 72468 66778 72480
rect 68278 72468 68284 72480
rect 66772 72440 68284 72468
rect 66772 72428 66778 72440
rect 68278 72428 68284 72440
rect 68336 72428 68342 72480
rect 106090 71856 106096 71868
rect 106016 71828 106096 71856
rect 106016 70780 106044 71828
rect 106090 71816 106096 71828
rect 106148 71816 106154 71868
rect 106182 71816 106188 71868
rect 106240 71816 106246 71868
rect 106090 71544 106096 71596
rect 106148 71584 106154 71596
rect 106200 71584 106228 71816
rect 107562 71748 107568 71800
rect 107620 71788 107626 71800
rect 167086 71788 167092 71800
rect 107620 71760 167092 71788
rect 107620 71748 107626 71760
rect 167086 71748 167092 71760
rect 167144 71748 167150 71800
rect 580166 71788 580172 71800
rect 202892 71760 580172 71788
rect 108482 71680 108488 71732
rect 108540 71720 108546 71732
rect 200298 71720 200304 71732
rect 108540 71692 200304 71720
rect 108540 71680 108546 71692
rect 200298 71680 200304 71692
rect 200356 71680 200362 71732
rect 201954 71680 201960 71732
rect 202012 71720 202018 71732
rect 202892 71720 202920 71760
rect 580166 71748 580172 71760
rect 580224 71748 580230 71800
rect 202012 71692 202920 71720
rect 202012 71680 202018 71692
rect 108574 71612 108580 71664
rect 108632 71652 108638 71664
rect 148962 71652 148968 71664
rect 108632 71624 148968 71652
rect 108632 71612 108638 71624
rect 148962 71612 148968 71624
rect 149020 71652 149026 71664
rect 200390 71652 200396 71664
rect 149020 71624 200396 71652
rect 149020 71612 149026 71624
rect 200390 71612 200396 71624
rect 200448 71612 200454 71664
rect 106148 71556 106228 71584
rect 106148 71544 106154 71556
rect 162854 71544 162860 71596
rect 162912 71584 162918 71596
rect 201494 71584 201500 71596
rect 162912 71556 201500 71584
rect 162912 71544 162918 71556
rect 201494 71544 201500 71556
rect 201552 71544 201558 71596
rect 164878 71476 164884 71528
rect 164936 71516 164942 71528
rect 201862 71516 201868 71528
rect 164936 71488 201868 71516
rect 164936 71476 164942 71488
rect 201862 71476 201868 71488
rect 201920 71476 201926 71528
rect 167454 71408 167460 71460
rect 167512 71448 167518 71460
rect 168006 71448 168012 71460
rect 167512 71420 168012 71448
rect 167512 71408 167518 71420
rect 168006 71408 168012 71420
rect 168064 71408 168070 71460
rect 200482 71340 200488 71392
rect 200540 71380 200546 71392
rect 201310 71380 201316 71392
rect 200540 71352 201316 71380
rect 200540 71340 200546 71352
rect 201310 71340 201316 71352
rect 201368 71340 201374 71392
rect 211890 71040 211896 71052
rect 209746 71012 211896 71040
rect 105998 70728 106004 70780
rect 106056 70728 106062 70780
rect 198826 70660 198832 70712
rect 198884 70700 198890 70712
rect 204806 70700 204812 70712
rect 198884 70672 204812 70700
rect 198884 70660 198890 70672
rect 204806 70660 204812 70672
rect 204864 70660 204870 70712
rect 198090 70592 198096 70644
rect 198148 70632 198154 70644
rect 209746 70632 209774 71012
rect 211890 71000 211896 71012
rect 211948 71000 211954 71052
rect 198148 70604 209774 70632
rect 198148 70592 198154 70604
rect 74534 70428 74540 70440
rect 74460 70400 74540 70428
rect 3602 70320 3608 70372
rect 3660 70360 3666 70372
rect 74460 70360 74488 70400
rect 74534 70388 74540 70400
rect 74592 70388 74598 70440
rect 75178 70388 75184 70440
rect 75236 70388 75242 70440
rect 76466 70388 76472 70440
rect 76524 70388 76530 70440
rect 87340 70400 87552 70428
rect 75196 70360 75224 70388
rect 3660 70332 74120 70360
rect 74460 70332 74534 70360
rect 3660 70320 3666 70332
rect 70394 70252 70400 70304
rect 70452 70292 70458 70304
rect 71268 70292 71274 70304
rect 70452 70264 71274 70292
rect 70452 70252 70458 70264
rect 71268 70252 71274 70264
rect 71326 70252 71332 70304
rect 71958 70252 71964 70304
rect 72016 70252 72022 70304
rect 72602 70252 72608 70304
rect 72660 70252 72666 70304
rect 73246 70252 73252 70304
rect 73304 70292 73310 70304
rect 73304 70264 73384 70292
rect 73304 70252 73310 70264
rect 71983 70156 72011 70252
rect 71976 70128 72011 70156
rect 67542 70048 67548 70100
rect 67600 70088 67606 70100
rect 70026 70088 70032 70100
rect 67600 70060 70032 70088
rect 67600 70048 67606 70060
rect 70026 70048 70032 70060
rect 70084 70048 70090 70100
rect 71976 69964 72004 70128
rect 72627 69964 72655 70252
rect 73356 69964 73384 70264
rect 73890 70252 73896 70304
rect 73948 70292 73954 70304
rect 73948 70264 74028 70292
rect 73948 70252 73954 70264
rect 74000 69964 74028 70264
rect 71958 69912 71964 69964
rect 72016 69912 72022 69964
rect 72602 69912 72608 69964
rect 72660 69912 72666 69964
rect 73338 69912 73344 69964
rect 73396 69912 73402 69964
rect 73982 69912 73988 69964
rect 74040 69912 74046 69964
rect 65978 69844 65984 69896
rect 66036 69884 66042 69896
rect 73706 69884 73712 69896
rect 66036 69856 73712 69884
rect 66036 69844 66042 69856
rect 73706 69844 73712 69856
rect 73764 69844 73770 69896
rect 74092 69884 74120 70332
rect 74506 70156 74534 70332
rect 75150 70332 75224 70360
rect 76484 70360 76512 70388
rect 76484 70332 76604 70360
rect 74506 70128 74580 70156
rect 74552 69964 74580 70128
rect 75150 69964 75178 70332
rect 76576 69964 76604 70332
rect 82866 70320 82872 70372
rect 82924 70320 82930 70372
rect 87340 70360 87368 70400
rect 84488 70332 87368 70360
rect 87524 70360 87552 70400
rect 87984 70400 88196 70428
rect 87984 70360 88012 70400
rect 87524 70332 88012 70360
rect 88168 70360 88196 70400
rect 97644 70400 97856 70428
rect 97644 70360 97672 70400
rect 88168 70332 97672 70360
rect 97828 70360 97856 70400
rect 99576 70400 99788 70428
rect 99576 70360 99604 70400
rect 97828 70332 99604 70360
rect 99760 70360 99788 70400
rect 100864 70400 101076 70428
rect 100864 70360 100892 70400
rect 101048 70394 101076 70400
rect 103164 70400 103468 70428
rect 99760 70332 100892 70360
rect 77110 70252 77116 70304
rect 77168 70252 77174 70304
rect 77754 70252 77760 70304
rect 77812 70252 77818 70304
rect 78398 70252 78404 70304
rect 78456 70252 78462 70304
rect 79042 70252 79048 70304
rect 79100 70252 79106 70304
rect 79686 70252 79692 70304
rect 79744 70252 79750 70304
rect 80330 70252 80336 70304
rect 80388 70252 80394 70304
rect 80974 70252 80980 70304
rect 81032 70252 81038 70304
rect 81618 70252 81624 70304
rect 81676 70252 81682 70304
rect 77135 70156 77163 70252
rect 77779 70156 77807 70252
rect 77128 70128 77163 70156
rect 77772 70128 77807 70156
rect 77128 69964 77156 70128
rect 77772 69964 77800 70128
rect 78423 69964 78451 70252
rect 79060 69964 79088 70252
rect 79704 69964 79732 70252
rect 80348 70224 80376 70252
rect 80992 70224 81020 70252
rect 81636 70224 81664 70252
rect 80348 70196 80468 70224
rect 80992 70196 81112 70224
rect 81636 70196 81756 70224
rect 80440 69964 80468 70196
rect 81084 69964 81112 70196
rect 81728 69964 81756 70196
rect 74534 69912 74540 69964
rect 74592 69912 74598 69964
rect 75150 69924 75184 69964
rect 75178 69912 75184 69924
rect 75236 69912 75242 69964
rect 76558 69912 76564 69964
rect 76616 69912 76622 69964
rect 77110 69912 77116 69964
rect 77168 69912 77174 69964
rect 77754 69912 77760 69964
rect 77812 69912 77818 69964
rect 78398 69912 78404 69964
rect 78456 69912 78462 69964
rect 79042 69912 79048 69964
rect 79100 69912 79106 69964
rect 79686 69912 79692 69964
rect 79744 69912 79750 69964
rect 80422 69912 80428 69964
rect 80480 69912 80486 69964
rect 81066 69912 81072 69964
rect 81124 69912 81130 69964
rect 81710 69912 81716 69964
rect 81768 69912 81774 69964
rect 82884 69924 82912 70320
rect 83550 70252 83556 70304
rect 83608 70252 83614 70304
rect 84194 70252 84200 70304
rect 84252 70252 84258 70304
rect 83568 70224 83596 70252
rect 83568 70196 83688 70224
rect 83660 69964 83688 70196
rect 84212 69964 84240 70252
rect 84488 70020 84516 70332
rect 100938 70320 100944 70372
rect 100996 70320 101002 70372
rect 101048 70366 101168 70394
rect 101140 70360 101168 70366
rect 101140 70332 102180 70360
rect 84854 70252 84860 70304
rect 84912 70252 84918 70304
rect 85482 70252 85488 70304
rect 85540 70252 85546 70304
rect 86126 70252 86132 70304
rect 86184 70252 86190 70304
rect 86770 70252 86776 70304
rect 86828 70252 86834 70304
rect 87414 70252 87420 70304
rect 87472 70252 87478 70304
rect 88058 70252 88064 70304
rect 88116 70252 88122 70304
rect 89346 70252 89352 70304
rect 89404 70252 89410 70304
rect 89990 70252 89996 70304
rect 90048 70252 90054 70304
rect 90634 70252 90640 70304
rect 90692 70252 90698 70304
rect 91278 70252 91284 70304
rect 91336 70252 91342 70304
rect 91922 70252 91928 70304
rect 91980 70252 91986 70304
rect 92566 70252 92572 70304
rect 92624 70252 92630 70304
rect 93210 70252 93216 70304
rect 93268 70252 93274 70304
rect 93854 70252 93860 70304
rect 93912 70252 93918 70304
rect 94514 70252 94520 70304
rect 94572 70252 94578 70304
rect 95786 70252 95792 70304
rect 95844 70252 95850 70304
rect 96430 70252 96436 70304
rect 96488 70252 96494 70304
rect 97074 70252 97080 70304
rect 97132 70252 97138 70304
rect 97718 70252 97724 70304
rect 97776 70252 97782 70304
rect 98362 70252 98368 70304
rect 98420 70252 98426 70304
rect 99006 70252 99012 70304
rect 99064 70252 99070 70304
rect 99650 70252 99656 70304
rect 99708 70252 99714 70304
rect 100294 70252 100300 70304
rect 100352 70252 100358 70304
rect 84872 70224 84900 70252
rect 84872 70196 84976 70224
rect 84304 69992 84516 70020
rect 82906 69912 82912 69924
rect 82964 69912 82970 69964
rect 83642 69912 83648 69964
rect 83700 69912 83706 69964
rect 84194 69912 84200 69964
rect 84252 69912 84258 69964
rect 84304 69884 84332 69992
rect 84948 69964 84976 70196
rect 85500 69964 85528 70252
rect 86144 69964 86172 70252
rect 86788 69964 86816 70252
rect 87432 69964 87460 70252
rect 88076 69964 88104 70252
rect 89364 69964 89392 70252
rect 84930 69912 84936 69964
rect 84988 69912 84994 69964
rect 85482 69912 85488 69964
rect 85540 69912 85546 69964
rect 86126 69912 86132 69964
rect 86184 69912 86190 69964
rect 86770 69912 86776 69964
rect 86828 69912 86834 69964
rect 87414 69912 87420 69964
rect 87472 69912 87478 69964
rect 88058 69912 88064 69964
rect 88116 69912 88122 69964
rect 89346 69912 89352 69964
rect 89404 69912 89410 69964
rect 90008 69896 90036 70252
rect 90652 69896 90680 70252
rect 91296 69896 91324 70252
rect 91940 69896 91968 70252
rect 92584 69896 92612 70252
rect 93228 69896 93256 70252
rect 93872 69896 93900 70252
rect 94532 70020 94560 70252
rect 94532 69992 94728 70020
rect 94700 69964 94728 69992
rect 95804 69964 95832 70252
rect 96448 69964 96476 70252
rect 97092 69964 97120 70252
rect 97736 69964 97764 70252
rect 98380 69964 98408 70252
rect 99024 69964 99052 70252
rect 99668 69964 99696 70252
rect 100312 69964 100340 70252
rect 100956 69964 100984 70320
rect 102152 69964 102180 70332
rect 102226 70252 102232 70304
rect 102284 70252 102290 70304
rect 102870 70252 102876 70304
rect 102928 70252 102934 70304
rect 102244 69964 102272 70252
rect 102888 69964 102916 70252
rect 103164 69964 103192 70400
rect 103440 70360 103468 70400
rect 166074 70388 166080 70440
rect 166132 70428 166138 70440
rect 168006 70428 168012 70440
rect 166132 70400 168012 70428
rect 166132 70388 166138 70400
rect 168006 70388 168012 70400
rect 168064 70388 168070 70440
rect 103440 70332 106320 70360
rect 103514 70252 103520 70304
rect 103572 70252 103578 70304
rect 104174 70252 104180 70304
rect 104232 70292 104238 70304
rect 104232 70264 104664 70292
rect 104232 70252 104238 70264
rect 103532 69964 103560 70252
rect 104636 69964 104664 70264
rect 104818 70252 104824 70304
rect 104876 70292 104882 70304
rect 104876 70264 105308 70292
rect 104876 70252 104882 70264
rect 105280 70156 105308 70264
rect 105462 70252 105468 70304
rect 105520 70292 105526 70304
rect 106182 70292 106188 70304
rect 105520 70264 106188 70292
rect 105520 70252 105526 70264
rect 106182 70252 106188 70264
rect 106240 70252 106246 70304
rect 106292 70292 106320 70332
rect 108022 70320 108028 70372
rect 108080 70360 108086 70372
rect 200114 70360 200120 70372
rect 108080 70332 200120 70360
rect 108080 70320 108086 70332
rect 200114 70320 200120 70332
rect 200172 70320 200178 70372
rect 106292 70264 161474 70292
rect 161446 70224 161474 70264
rect 164786 70252 164792 70304
rect 164844 70292 164850 70304
rect 204438 70292 204444 70304
rect 164844 70264 204444 70292
rect 164844 70252 164850 70264
rect 204438 70252 204444 70264
rect 204496 70252 204502 70304
rect 165154 70224 165160 70236
rect 161446 70196 165160 70224
rect 165154 70184 165160 70196
rect 165212 70184 165218 70236
rect 165246 70184 165252 70236
rect 165304 70224 165310 70236
rect 203242 70224 203248 70236
rect 165304 70196 203248 70224
rect 165304 70184 165310 70196
rect 203242 70184 203248 70196
rect 203300 70184 203306 70236
rect 110322 70156 110328 70168
rect 105280 70128 110328 70156
rect 110322 70116 110328 70128
rect 110380 70156 110386 70168
rect 200390 70156 200396 70168
rect 110380 70128 200396 70156
rect 110380 70116 110386 70128
rect 200390 70116 200396 70128
rect 200448 70116 200454 70168
rect 108666 70048 108672 70100
rect 108724 70088 108730 70100
rect 200022 70088 200028 70100
rect 108724 70060 200028 70088
rect 108724 70048 108730 70060
rect 200022 70048 200028 70060
rect 200080 70048 200086 70100
rect 115750 69980 115756 70032
rect 115808 70020 115814 70032
rect 200482 70020 200488 70032
rect 115808 69992 200488 70020
rect 115808 69980 115814 69992
rect 200482 69980 200488 69992
rect 200540 69980 200546 70032
rect 94682 69912 94688 69964
rect 94740 69912 94746 69964
rect 95786 69912 95792 69964
rect 95844 69912 95850 69964
rect 96430 69912 96436 69964
rect 96488 69912 96494 69964
rect 97074 69912 97080 69964
rect 97132 69912 97138 69964
rect 97718 69912 97724 69964
rect 97776 69912 97782 69964
rect 98362 69912 98368 69964
rect 98420 69912 98426 69964
rect 99006 69912 99012 69964
rect 99064 69912 99070 69964
rect 99650 69912 99656 69964
rect 99708 69912 99714 69964
rect 100294 69912 100300 69964
rect 100352 69912 100358 69964
rect 100938 69912 100944 69964
rect 100996 69912 101002 69964
rect 102134 69912 102140 69964
rect 102192 69912 102198 69964
rect 102226 69912 102232 69964
rect 102284 69912 102290 69964
rect 102870 69912 102876 69964
rect 102928 69912 102934 69964
rect 103146 69912 103152 69964
rect 103204 69912 103210 69964
rect 103514 69912 103520 69964
rect 103572 69912 103578 69964
rect 104618 69912 104624 69964
rect 104676 69912 104682 69964
rect 165062 69912 165068 69964
rect 165120 69952 165126 69964
rect 201770 69952 201776 69964
rect 165120 69924 201776 69952
rect 165120 69912 165126 69924
rect 201770 69912 201776 69924
rect 201828 69912 201834 69964
rect 74092 69856 84332 69884
rect 84470 69844 84476 69896
rect 84528 69884 84534 69896
rect 89898 69884 89904 69896
rect 84528 69856 89904 69884
rect 84528 69844 84534 69856
rect 89898 69844 89904 69856
rect 89956 69844 89962 69896
rect 89990 69844 89996 69896
rect 90048 69844 90054 69896
rect 90634 69844 90640 69896
rect 90692 69844 90698 69896
rect 91278 69844 91284 69896
rect 91336 69844 91342 69896
rect 91922 69844 91928 69896
rect 91980 69844 91986 69896
rect 92566 69844 92572 69896
rect 92624 69844 92630 69896
rect 93210 69844 93216 69896
rect 93268 69844 93274 69896
rect 93854 69844 93860 69896
rect 93912 69844 93918 69896
rect 165522 69884 165528 69896
rect 94424 69856 165528 69884
rect 70302 69776 70308 69828
rect 70360 69816 70366 69828
rect 75362 69816 75368 69828
rect 70360 69788 75368 69816
rect 70360 69776 70366 69788
rect 75362 69776 75368 69788
rect 75420 69776 75426 69828
rect 84010 69776 84016 69828
rect 84068 69816 84074 69828
rect 84068 69788 89714 69816
rect 84068 69776 84074 69788
rect 68554 69708 68560 69760
rect 68612 69748 68618 69760
rect 68612 69720 75224 69748
rect 68612 69708 68618 69720
rect 68370 69640 68376 69692
rect 68428 69680 68434 69692
rect 75196 69680 75224 69720
rect 75270 69708 75276 69760
rect 75328 69748 75334 69760
rect 89686 69748 89714 69788
rect 94424 69748 94452 69856
rect 165522 69844 165528 69856
rect 165580 69844 165586 69896
rect 166718 69844 166724 69896
rect 166776 69884 166782 69896
rect 195238 69884 195244 69896
rect 166776 69856 195244 69884
rect 166776 69844 166782 69856
rect 195238 69844 195244 69856
rect 195296 69844 195302 69896
rect 201678 69884 201684 69896
rect 195348 69856 201684 69884
rect 107286 69816 107292 69828
rect 75328 69720 84240 69748
rect 89686 69720 94452 69748
rect 94516 69788 107292 69816
rect 75328 69708 75334 69720
rect 84212 69680 84240 69720
rect 94516 69680 94544 69788
rect 107286 69776 107292 69788
rect 107344 69776 107350 69828
rect 166534 69776 166540 69828
rect 166592 69816 166598 69828
rect 195348 69816 195376 69856
rect 201678 69844 201684 69856
rect 201736 69844 201742 69896
rect 166592 69788 195376 69816
rect 166592 69776 166598 69788
rect 195422 69776 195428 69828
rect 195480 69816 195486 69828
rect 202230 69816 202236 69828
rect 195480 69788 202236 69816
rect 195480 69776 195486 69788
rect 202230 69776 202236 69788
rect 202288 69776 202294 69828
rect 102134 69708 102140 69760
rect 102192 69748 102198 69760
rect 106458 69748 106464 69760
rect 102192 69720 106464 69748
rect 102192 69708 102198 69720
rect 106458 69708 106464 69720
rect 106516 69708 106522 69760
rect 166442 69708 166448 69760
rect 166500 69748 166506 69760
rect 201586 69748 201592 69760
rect 166500 69720 201592 69748
rect 166500 69708 166506 69720
rect 201586 69708 201592 69720
rect 201644 69708 201650 69760
rect 68428 69652 70394 69680
rect 75196 69652 84148 69680
rect 84212 69652 94544 69680
rect 68428 69640 68434 69652
rect 70366 69612 70394 69652
rect 75270 69612 75276 69624
rect 70366 69584 75276 69612
rect 75270 69572 75276 69584
rect 75328 69572 75334 69624
rect 75362 69572 75368 69624
rect 75420 69612 75426 69624
rect 84010 69612 84016 69624
rect 75420 69584 84016 69612
rect 75420 69572 75426 69584
rect 84010 69572 84016 69584
rect 84068 69572 84074 69624
rect 84120 69612 84148 69652
rect 166902 69640 166908 69692
rect 166960 69680 166966 69692
rect 202138 69680 202144 69692
rect 166960 69652 202144 69680
rect 166960 69640 166966 69652
rect 202138 69640 202144 69652
rect 202196 69640 202202 69692
rect 202782 69640 202788 69692
rect 202840 69680 202846 69692
rect 210602 69680 210608 69692
rect 202840 69652 210608 69680
rect 202840 69640 202846 69652
rect 210602 69640 210608 69652
rect 210660 69640 210666 69692
rect 84120 69584 89714 69612
rect 73706 69504 73712 69556
rect 73764 69544 73770 69556
rect 84470 69544 84476 69556
rect 73764 69516 84476 69544
rect 73764 69504 73770 69516
rect 84470 69504 84476 69516
rect 84528 69504 84534 69556
rect 89686 69544 89714 69584
rect 89898 69572 89904 69624
rect 89956 69612 89962 69624
rect 103146 69612 103152 69624
rect 89956 69584 103152 69612
rect 89956 69572 89962 69584
rect 103146 69572 103152 69584
rect 103204 69572 103210 69624
rect 166626 69572 166632 69624
rect 166684 69612 166690 69624
rect 166684 69584 180794 69612
rect 166684 69572 166690 69584
rect 107102 69544 107108 69556
rect 89686 69516 107108 69544
rect 107102 69504 107108 69516
rect 107160 69504 107166 69556
rect 180766 69544 180794 69584
rect 202414 69544 202420 69556
rect 180766 69516 202420 69544
rect 202414 69504 202420 69516
rect 202472 69504 202478 69556
rect 202690 69436 202696 69488
rect 202748 69476 202754 69488
rect 206094 69476 206100 69488
rect 202748 69448 206100 69476
rect 202748 69436 202754 69448
rect 206094 69436 206100 69448
rect 206152 69436 206158 69488
rect 104618 69096 104624 69148
rect 104676 69136 104682 69148
rect 113174 69136 113180 69148
rect 104676 69108 113180 69136
rect 104676 69096 104682 69108
rect 113174 69096 113180 69108
rect 113232 69136 113238 69148
rect 113542 69136 113548 69148
rect 113232 69108 113548 69136
rect 113232 69096 113238 69108
rect 113542 69096 113548 69108
rect 113600 69096 113606 69148
rect 106182 69028 106188 69080
rect 106240 69068 106246 69080
rect 115750 69068 115756 69080
rect 106240 69040 115756 69068
rect 106240 69028 106246 69040
rect 115750 69028 115756 69040
rect 115808 69028 115814 69080
rect 166258 69028 166264 69080
rect 166316 69068 166322 69080
rect 178034 69068 178040 69080
rect 166316 69040 178040 69068
rect 166316 69028 166322 69040
rect 178034 69028 178040 69040
rect 178092 69068 178098 69080
rect 179046 69068 179052 69080
rect 178092 69040 179052 69068
rect 178092 69028 178098 69040
rect 179046 69028 179052 69040
rect 179104 69028 179110 69080
rect 97718 68960 97724 69012
rect 97776 69000 97782 69012
rect 104158 69000 104164 69012
rect 97776 68972 104164 69000
rect 97776 68960 97782 68972
rect 104158 68960 104164 68972
rect 104216 68960 104222 69012
rect 163958 69000 163964 69012
rect 161446 68972 163964 69000
rect 63218 68892 63224 68944
rect 63276 68932 63282 68944
rect 71958 68932 71964 68944
rect 63276 68904 71964 68932
rect 63276 68892 63282 68904
rect 71958 68892 71964 68904
rect 72016 68932 72022 68944
rect 161446 68932 161474 68972
rect 163958 68960 163964 68972
rect 164016 69000 164022 69012
rect 171778 69000 171784 69012
rect 164016 68972 171784 69000
rect 164016 68960 164022 68972
rect 171778 68960 171784 68972
rect 171836 68960 171842 69012
rect 196618 68960 196624 69012
rect 196676 69000 196682 69012
rect 202782 69000 202788 69012
rect 196676 68972 202788 69000
rect 196676 68960 196682 68972
rect 202782 68960 202788 68972
rect 202840 68960 202846 69012
rect 212534 69000 212540 69012
rect 209746 68972 212540 69000
rect 72016 68904 161474 68932
rect 72016 68892 72022 68904
rect 166258 68892 166264 68944
rect 166316 68932 166322 68944
rect 184198 68932 184204 68944
rect 166316 68904 184204 68932
rect 166316 68892 166322 68904
rect 184198 68892 184204 68904
rect 184256 68892 184262 68944
rect 192570 68892 192576 68944
rect 192628 68932 192634 68944
rect 202598 68932 202604 68944
rect 192628 68904 202604 68932
rect 192628 68892 192634 68904
rect 202598 68892 202604 68904
rect 202656 68892 202662 68944
rect 61838 68824 61844 68876
rect 61896 68864 61902 68876
rect 77754 68864 77760 68876
rect 61896 68836 77760 68864
rect 61896 68824 61902 68836
rect 77754 68824 77760 68836
rect 77812 68824 77818 68876
rect 91922 68824 91928 68876
rect 91980 68864 91986 68876
rect 95142 68864 95148 68876
rect 91980 68836 95148 68864
rect 91980 68824 91986 68836
rect 95142 68824 95148 68836
rect 95200 68824 95206 68876
rect 97074 68824 97080 68876
rect 97132 68864 97138 68876
rect 109126 68864 109132 68876
rect 97132 68836 109132 68864
rect 97132 68824 97138 68836
rect 109126 68824 109132 68836
rect 109184 68864 109190 68876
rect 209746 68864 209774 68972
rect 212534 68960 212540 68972
rect 212592 69000 212598 69012
rect 213822 69000 213828 69012
rect 212592 68972 213828 69000
rect 212592 68960 212598 68972
rect 213822 68960 213828 68972
rect 213880 68960 213886 69012
rect 109184 68836 196204 68864
rect 109184 68824 109190 68836
rect 92566 68756 92572 68808
rect 92624 68796 92630 68808
rect 106274 68796 106280 68808
rect 92624 68768 106280 68796
rect 92624 68756 92630 68768
rect 106274 68756 106280 68768
rect 106332 68796 106338 68808
rect 193214 68796 193220 68808
rect 106332 68768 193220 68796
rect 106332 68756 106338 68768
rect 193214 68756 193220 68768
rect 193272 68756 193278 68808
rect 196176 68796 196204 68836
rect 198752 68836 209774 68864
rect 197722 68796 197728 68808
rect 196176 68768 197728 68796
rect 197722 68756 197728 68768
rect 197780 68796 197786 68808
rect 198642 68796 198648 68808
rect 197780 68768 198648 68796
rect 197780 68756 197786 68768
rect 198642 68756 198648 68768
rect 198700 68756 198706 68808
rect 65794 68688 65800 68740
rect 65852 68728 65858 68740
rect 77110 68728 77116 68740
rect 65852 68700 77116 68728
rect 65852 68688 65858 68700
rect 77110 68688 77116 68700
rect 77168 68728 77174 68740
rect 163774 68728 163780 68740
rect 77168 68700 163780 68728
rect 77168 68688 77174 68700
rect 163774 68688 163780 68700
rect 163832 68728 163838 68740
rect 177390 68728 177396 68740
rect 163832 68700 177396 68728
rect 163832 68688 163838 68700
rect 177390 68688 177396 68700
rect 177448 68688 177454 68740
rect 198366 68728 198372 68740
rect 180766 68700 198372 68728
rect 76558 68620 76564 68672
rect 76616 68660 76622 68672
rect 104066 68660 104072 68672
rect 76616 68632 104072 68660
rect 76616 68620 76622 68632
rect 104066 68620 104072 68632
rect 104124 68620 104130 68672
rect 104158 68620 104164 68672
rect 104216 68660 104222 68672
rect 113266 68660 113272 68672
rect 104216 68632 113272 68660
rect 104216 68620 104222 68632
rect 113266 68620 113272 68632
rect 113324 68660 113330 68672
rect 180766 68660 180794 68700
rect 198366 68688 198372 68700
rect 198424 68728 198430 68740
rect 198752 68728 198780 68836
rect 198424 68700 198780 68728
rect 198424 68688 198430 68700
rect 113324 68632 180794 68660
rect 113324 68620 113330 68632
rect 193858 68620 193864 68672
rect 193916 68660 193922 68672
rect 194410 68660 194416 68672
rect 193916 68632 194416 68660
rect 193916 68620 193922 68632
rect 194410 68620 194416 68632
rect 194468 68660 194474 68672
rect 202690 68660 202696 68672
rect 194468 68632 202696 68660
rect 194468 68620 194474 68632
rect 202690 68620 202696 68632
rect 202748 68620 202754 68672
rect 93210 68552 93216 68604
rect 93268 68592 93274 68604
rect 110598 68592 110604 68604
rect 93268 68564 110604 68592
rect 93268 68552 93274 68564
rect 110598 68552 110604 68564
rect 110656 68592 110662 68604
rect 193876 68592 193904 68620
rect 110656 68564 193904 68592
rect 110656 68552 110662 68564
rect 81066 68484 81072 68536
rect 81124 68524 81130 68536
rect 156690 68524 156696 68536
rect 81124 68496 156696 68524
rect 81124 68484 81130 68496
rect 156690 68484 156696 68496
rect 156748 68524 156754 68536
rect 181438 68524 181444 68536
rect 156748 68496 181444 68524
rect 156748 68484 156754 68496
rect 181438 68484 181444 68496
rect 181496 68484 181502 68536
rect 193214 68484 193220 68536
rect 193272 68524 193278 68536
rect 194318 68524 194324 68536
rect 193272 68496 194324 68524
rect 193272 68484 193278 68496
rect 194318 68484 194324 68496
rect 194376 68524 194382 68536
rect 198826 68524 198832 68536
rect 194376 68496 198832 68524
rect 194376 68484 194382 68496
rect 198826 68484 198832 68496
rect 198884 68484 198890 68536
rect 86770 68416 86776 68468
rect 86828 68456 86834 68468
rect 111794 68456 111800 68468
rect 86828 68428 111800 68456
rect 86828 68416 86834 68428
rect 111794 68416 111800 68428
rect 111852 68456 111858 68468
rect 187418 68456 187424 68468
rect 111852 68428 187424 68456
rect 111852 68416 111858 68428
rect 187418 68416 187424 68428
rect 187476 68416 187482 68468
rect 72602 68348 72608 68400
rect 72660 68388 72666 68400
rect 108114 68388 108120 68400
rect 72660 68360 108120 68388
rect 72660 68348 72666 68360
rect 108114 68348 108120 68360
rect 108172 68388 108178 68400
rect 172974 68388 172980 68400
rect 108172 68360 172980 68388
rect 108172 68348 108178 68360
rect 172974 68348 172980 68360
rect 173032 68348 173038 68400
rect 213822 68348 213828 68400
rect 213880 68388 213886 68400
rect 293954 68388 293960 68400
rect 213880 68360 293960 68388
rect 213880 68348 213886 68360
rect 293954 68348 293960 68360
rect 294012 68348 294018 68400
rect 96430 68280 96436 68332
rect 96488 68320 96494 68332
rect 104158 68320 104164 68332
rect 96488 68292 104164 68320
rect 96488 68280 96494 68292
rect 104158 68280 104164 68292
rect 104216 68280 104222 68332
rect 104250 68280 104256 68332
rect 104308 68320 104314 68332
rect 112438 68320 112444 68332
rect 104308 68292 112444 68320
rect 104308 68280 104314 68292
rect 112438 68280 112444 68292
rect 112496 68320 112502 68332
rect 175918 68320 175924 68332
rect 112496 68292 175924 68320
rect 112496 68280 112502 68292
rect 175918 68280 175924 68292
rect 175976 68280 175982 68332
rect 202598 68280 202604 68332
rect 202656 68320 202662 68332
rect 204162 68320 204168 68332
rect 202656 68292 204168 68320
rect 202656 68280 202662 68292
rect 204162 68280 204168 68292
rect 204220 68320 204226 68332
rect 350534 68320 350540 68332
rect 204220 68292 350540 68320
rect 204220 68280 204226 68292
rect 350534 68280 350540 68292
rect 350592 68280 350598 68332
rect 86126 68212 86132 68264
rect 86184 68252 86190 68264
rect 123570 68252 123576 68264
rect 86184 68224 123576 68252
rect 86184 68212 86190 68224
rect 123570 68212 123576 68224
rect 123628 68252 123634 68264
rect 186958 68252 186964 68264
rect 123628 68224 186964 68252
rect 123628 68212 123634 68224
rect 186958 68212 186964 68224
rect 187016 68212 187022 68264
rect 188338 68184 188344 68196
rect 132466 68156 188344 68184
rect 87414 68076 87420 68128
rect 87472 68116 87478 68128
rect 127802 68116 127808 68128
rect 87472 68088 127808 68116
rect 87472 68076 87478 68088
rect 127802 68076 127808 68088
rect 127860 68116 127866 68128
rect 132466 68116 132494 68156
rect 188338 68144 188344 68156
rect 188396 68144 188402 68196
rect 127860 68088 132494 68116
rect 127860 68076 127866 68088
rect 70486 68008 70492 68060
rect 70544 68048 70550 68060
rect 170490 68048 170496 68060
rect 70544 68020 170496 68048
rect 70544 68008 70550 68020
rect 170490 68008 170496 68020
rect 170548 68048 170554 68060
rect 170674 68048 170680 68060
rect 170548 68020 170680 68048
rect 170548 68008 170554 68020
rect 170674 68008 170680 68020
rect 170732 68008 170738 68060
rect 104158 67940 104164 67992
rect 104216 67980 104222 67992
rect 110506 67980 110512 67992
rect 104216 67952 110512 67980
rect 104216 67940 104222 67952
rect 110506 67940 110512 67952
rect 110564 67940 110570 67992
rect 105998 67572 106004 67584
rect 99346 67544 106004 67572
rect 68830 67328 68836 67380
rect 68888 67368 68894 67380
rect 99346 67368 99374 67544
rect 105998 67532 106004 67544
rect 106056 67532 106062 67584
rect 113082 67532 113088 67584
rect 113140 67572 113146 67584
rect 200666 67572 200672 67584
rect 113140 67544 200672 67572
rect 113140 67532 113146 67544
rect 200666 67532 200672 67544
rect 200724 67532 200730 67584
rect 204438 67532 204444 67584
rect 204496 67572 204502 67584
rect 233878 67572 233884 67584
rect 204496 67544 233884 67572
rect 204496 67532 204502 67544
rect 233878 67532 233884 67544
rect 233936 67532 233942 67584
rect 99650 67464 99656 67516
rect 99708 67504 99714 67516
rect 110414 67504 110420 67516
rect 99708 67476 110420 67504
rect 99708 67464 99714 67476
rect 110414 67464 110420 67476
rect 110472 67504 110478 67516
rect 199378 67504 199384 67516
rect 110472 67476 199384 67504
rect 110472 67464 110478 67476
rect 199378 67464 199384 67476
rect 199436 67504 199442 67516
rect 215294 67504 215300 67516
rect 199436 67476 215300 67504
rect 199436 67464 199442 67476
rect 215294 67464 215300 67476
rect 215352 67464 215358 67516
rect 102870 67396 102876 67448
rect 102928 67436 102934 67448
rect 102928 67408 122834 67436
rect 102928 67396 102934 67408
rect 115198 67368 115204 67380
rect 68888 67340 99374 67368
rect 104084 67340 115204 67368
rect 68888 67328 68894 67340
rect 2866 67260 2872 67312
rect 2924 67300 2930 67312
rect 103974 67300 103980 67312
rect 2924 67272 103980 67300
rect 2924 67260 2930 67272
rect 103974 67260 103980 67272
rect 104032 67260 104038 67312
rect 80422 67192 80428 67244
rect 80480 67232 80486 67244
rect 104084 67232 104112 67340
rect 115198 67328 115204 67340
rect 115256 67368 115262 67380
rect 115842 67368 115848 67380
rect 115256 67340 115848 67368
rect 115256 67328 115262 67340
rect 115842 67328 115848 67340
rect 115900 67328 115906 67380
rect 122806 67368 122834 67408
rect 175826 67396 175832 67448
rect 175884 67436 175890 67448
rect 258718 67436 258724 67448
rect 175884 67408 258724 67436
rect 175884 67396 175890 67408
rect 258718 67396 258724 67408
rect 258776 67396 258782 67448
rect 123754 67368 123760 67380
rect 122806 67340 123760 67368
rect 123754 67328 123760 67340
rect 123812 67368 123818 67380
rect 200574 67368 200580 67380
rect 123812 67340 200580 67368
rect 123812 67328 123818 67340
rect 200574 67328 200580 67340
rect 200632 67328 200638 67380
rect 104158 67260 104164 67312
rect 104216 67300 104222 67312
rect 106550 67300 106556 67312
rect 104216 67272 106556 67300
rect 104216 67260 104222 67272
rect 106550 67260 106556 67272
rect 106608 67260 106614 67312
rect 109034 67300 109040 67312
rect 108947 67272 109040 67300
rect 109006 67260 109040 67272
rect 109092 67300 109098 67312
rect 182910 67300 182916 67312
rect 109092 67272 182916 67300
rect 109092 67260 109098 67272
rect 182910 67260 182916 67272
rect 182968 67300 182974 67312
rect 204438 67300 204444 67312
rect 182968 67272 204444 67300
rect 182968 67260 182974 67272
rect 204438 67260 204444 67272
rect 204496 67260 204502 67312
rect 109006 67232 109034 67260
rect 80480 67204 104112 67232
rect 104176 67204 109034 67232
rect 80480 67192 80486 67204
rect 82906 67124 82912 67176
rect 82964 67164 82970 67176
rect 104176 67164 104204 67204
rect 127618 67192 127624 67244
rect 127676 67232 127682 67244
rect 199010 67232 199016 67244
rect 127676 67204 199016 67232
rect 127676 67192 127682 67204
rect 199010 67192 199016 67204
rect 199068 67192 199074 67244
rect 82964 67136 104204 67164
rect 82964 67124 82970 67136
rect 109034 67124 109040 67176
rect 109092 67164 109098 67176
rect 109678 67164 109684 67176
rect 109092 67136 109684 67164
rect 109092 67124 109098 67136
rect 109678 67124 109684 67136
rect 109736 67164 109742 67176
rect 173894 67164 173900 67176
rect 109736 67136 173900 67164
rect 109736 67124 109742 67136
rect 173894 67124 173900 67136
rect 173952 67124 173958 67176
rect 187418 67124 187424 67176
rect 187476 67164 187482 67176
rect 203426 67164 203432 67176
rect 187476 67136 203432 67164
rect 187476 67124 187482 67136
rect 203426 67124 203432 67136
rect 203484 67124 203490 67176
rect 95786 67056 95792 67108
rect 95844 67096 95850 67108
rect 131758 67096 131764 67108
rect 95844 67068 131764 67096
rect 95844 67056 95850 67068
rect 131758 67056 131764 67068
rect 131816 67096 131822 67108
rect 196434 67096 196440 67108
rect 131816 67068 196440 67096
rect 131816 67056 131822 67068
rect 196434 67056 196440 67068
rect 196492 67056 196498 67108
rect 93854 66988 93860 67040
rect 93912 67028 93918 67040
rect 130378 67028 130384 67040
rect 93912 67000 130384 67028
rect 93912 66988 93918 67000
rect 130378 66988 130384 67000
rect 130436 67028 130442 67040
rect 194502 67028 194508 67040
rect 130436 67000 194508 67028
rect 130436 66988 130442 67000
rect 194502 66988 194508 67000
rect 194560 66988 194566 67040
rect 99006 66920 99012 66972
rect 99064 66960 99070 66972
rect 137278 66960 137284 66972
rect 99064 66932 137284 66960
rect 99064 66920 99070 66932
rect 137278 66920 137284 66932
rect 137336 66960 137342 66972
rect 199654 66960 199660 66972
rect 137336 66932 199660 66960
rect 137336 66920 137342 66932
rect 199654 66920 199660 66932
rect 199712 66920 199718 66972
rect 100294 66852 100300 66904
rect 100352 66892 100358 66904
rect 142982 66892 142988 66904
rect 100352 66864 142988 66892
rect 100352 66852 100358 66864
rect 142982 66852 142988 66864
rect 143040 66892 143046 66904
rect 198734 66892 198740 66904
rect 143040 66864 198740 66892
rect 143040 66852 143046 66864
rect 198734 66852 198740 66864
rect 198792 66852 198798 66904
rect 215294 66852 215300 66904
rect 215352 66892 215358 66904
rect 216398 66892 216404 66904
rect 215352 66864 216404 66892
rect 215352 66852 215358 66864
rect 216398 66852 216404 66864
rect 216456 66892 216462 66904
rect 349246 66892 349252 66904
rect 216456 66864 349252 66892
rect 216456 66852 216462 66864
rect 349246 66852 349252 66864
rect 349304 66852 349310 66904
rect 98362 66784 98368 66836
rect 98420 66824 98426 66836
rect 127618 66824 127624 66836
rect 98420 66796 127624 66824
rect 98420 66784 98426 66796
rect 127618 66784 127624 66796
rect 127676 66784 127682 66836
rect 165430 66784 165436 66836
rect 165488 66824 165494 66836
rect 185578 66824 185584 66836
rect 165488 66796 185584 66824
rect 165488 66784 165494 66796
rect 185578 66784 185584 66796
rect 185636 66784 185642 66836
rect 67818 66716 67824 66768
rect 67876 66756 67882 66768
rect 107378 66756 107384 66768
rect 67876 66728 107384 66756
rect 67876 66716 67882 66728
rect 107378 66716 107384 66728
rect 107436 66716 107442 66768
rect 115842 66716 115848 66768
rect 115900 66756 115906 66768
rect 180978 66756 180984 66768
rect 115900 66728 180984 66756
rect 115900 66716 115906 66728
rect 180978 66716 180984 66728
rect 181036 66716 181042 66768
rect 68922 66648 68928 66700
rect 68980 66688 68986 66700
rect 106090 66688 106096 66700
rect 68980 66660 106096 66688
rect 68980 66648 68986 66660
rect 106090 66648 106096 66660
rect 106148 66648 106154 66700
rect 73982 66580 73988 66632
rect 74040 66620 74046 66632
rect 109034 66620 109040 66632
rect 74040 66592 109040 66620
rect 74040 66580 74046 66592
rect 109034 66580 109040 66592
rect 109092 66580 109098 66632
rect 85482 66172 85488 66224
rect 85540 66212 85546 66224
rect 108390 66212 108396 66224
rect 85540 66184 108396 66212
rect 85540 66172 85546 66184
rect 108390 66172 108396 66184
rect 108448 66172 108454 66224
rect 162118 66172 162124 66224
rect 162176 66212 162182 66224
rect 208394 66212 208400 66224
rect 162176 66184 208400 66212
rect 162176 66172 162182 66184
rect 208394 66172 208400 66184
rect 208452 66172 208458 66224
rect 91278 66104 91284 66156
rect 91336 66144 91342 66156
rect 123662 66144 123668 66156
rect 91336 66116 123668 66144
rect 91336 66104 91342 66116
rect 123662 66104 123668 66116
rect 123720 66144 123726 66156
rect 191926 66144 191932 66156
rect 123720 66116 191932 66144
rect 123720 66104 123726 66116
rect 191926 66104 191932 66116
rect 191984 66104 191990 66156
rect 83642 66036 83648 66088
rect 83700 66076 83706 66088
rect 121454 66076 121460 66088
rect 83700 66048 121460 66076
rect 83700 66036 83706 66048
rect 121454 66036 121460 66048
rect 121512 66036 121518 66088
rect 125318 66036 125324 66088
rect 125376 66076 125382 66088
rect 125502 66076 125508 66088
rect 125376 66048 125508 66076
rect 125376 66036 125382 66048
rect 125502 66036 125508 66048
rect 125560 66076 125566 66088
rect 191098 66076 191104 66088
rect 125560 66048 191104 66076
rect 125560 66036 125566 66048
rect 191098 66036 191104 66048
rect 191156 66076 191162 66088
rect 191282 66076 191288 66088
rect 191156 66048 191288 66076
rect 191156 66036 191162 66048
rect 191282 66036 191288 66048
rect 191340 66036 191346 66088
rect 94682 65968 94688 66020
rect 94740 66008 94746 66020
rect 133322 66008 133328 66020
rect 94740 65980 133328 66008
rect 94740 65968 94746 65980
rect 133322 65968 133328 65980
rect 133380 66008 133386 66020
rect 133782 66008 133788 66020
rect 133380 65980 133788 66008
rect 133380 65968 133386 65980
rect 133782 65968 133788 65980
rect 133840 65968 133846 66020
rect 135162 65968 135168 66020
rect 135220 66008 135226 66020
rect 200758 66008 200764 66020
rect 135220 65980 200764 66008
rect 135220 65968 135226 65980
rect 200758 65968 200764 65980
rect 200816 65968 200822 66020
rect 67910 65900 67916 65952
rect 67968 65940 67974 65952
rect 107194 65940 107200 65952
rect 67968 65912 107200 65940
rect 67968 65900 67974 65912
rect 107194 65900 107200 65912
rect 107252 65900 107258 65952
rect 162302 65900 162308 65952
rect 162360 65940 162366 65952
rect 203150 65940 203156 65952
rect 162360 65912 203156 65940
rect 162360 65900 162366 65912
rect 203150 65900 203156 65912
rect 203208 65900 203214 65952
rect 84930 65832 84936 65884
rect 84988 65872 84994 65884
rect 123478 65872 123484 65884
rect 84988 65844 123484 65872
rect 84988 65832 84994 65844
rect 123478 65832 123484 65844
rect 123536 65872 123542 65884
rect 124122 65872 124128 65884
rect 123536 65844 124128 65872
rect 123536 65832 123542 65844
rect 124122 65832 124128 65844
rect 124180 65832 124186 65884
rect 126882 65832 126888 65884
rect 126940 65872 126946 65884
rect 189994 65872 190000 65884
rect 126940 65844 190000 65872
rect 126940 65832 126946 65844
rect 189994 65832 190000 65844
rect 190052 65832 190058 65884
rect 75178 65764 75184 65816
rect 75236 65804 75242 65816
rect 110874 65804 110880 65816
rect 75236 65776 110880 65804
rect 75236 65764 75242 65776
rect 110874 65764 110880 65776
rect 110932 65804 110938 65816
rect 111150 65804 111156 65816
rect 110932 65776 111156 65804
rect 110932 65764 110938 65776
rect 111150 65764 111156 65776
rect 111208 65764 111214 65816
rect 121454 65764 121460 65816
rect 121512 65804 121518 65816
rect 122098 65804 122104 65816
rect 121512 65776 122104 65804
rect 121512 65764 121518 65776
rect 122098 65764 122104 65776
rect 122156 65804 122162 65816
rect 183554 65804 183560 65816
rect 122156 65776 183560 65804
rect 122156 65764 122162 65776
rect 183554 65764 183560 65776
rect 183612 65764 183618 65816
rect 89990 65696 89996 65748
rect 90048 65736 90054 65748
rect 126330 65736 126336 65748
rect 90048 65708 126336 65736
rect 90048 65696 90054 65708
rect 126330 65696 126336 65708
rect 126388 65736 126394 65748
rect 126882 65736 126888 65748
rect 126388 65708 126888 65736
rect 126388 65696 126394 65708
rect 126882 65696 126888 65708
rect 126940 65696 126946 65748
rect 133782 65696 133788 65748
rect 133840 65736 133846 65748
rect 195146 65736 195152 65748
rect 133840 65708 195152 65736
rect 133840 65696 133846 65708
rect 195146 65696 195152 65708
rect 195204 65696 195210 65748
rect 208394 65696 208400 65748
rect 208452 65736 208458 65748
rect 209038 65736 209044 65748
rect 208452 65708 209044 65736
rect 208452 65696 208458 65708
rect 209038 65696 209044 65708
rect 209096 65696 209102 65748
rect 124122 65628 124128 65680
rect 124180 65668 124186 65680
rect 184842 65668 184848 65680
rect 124180 65640 184848 65668
rect 124180 65628 124186 65640
rect 184842 65628 184848 65640
rect 184900 65628 184906 65680
rect 102226 65560 102232 65612
rect 102284 65600 102290 65612
rect 134702 65600 134708 65612
rect 102284 65572 134708 65600
rect 102284 65560 102290 65572
rect 134702 65560 134708 65572
rect 134760 65600 134766 65612
rect 135162 65600 135168 65612
rect 134760 65572 135168 65600
rect 134760 65560 134766 65572
rect 135162 65560 135168 65572
rect 135220 65560 135226 65612
rect 162394 65560 162400 65612
rect 162452 65600 162458 65612
rect 203334 65600 203340 65612
rect 162452 65572 203340 65600
rect 162452 65560 162458 65572
rect 203334 65560 203340 65572
rect 203392 65560 203398 65612
rect 79042 65492 79048 65544
rect 79100 65532 79106 65544
rect 107930 65532 107936 65544
rect 79100 65504 107936 65532
rect 79100 65492 79106 65504
rect 107930 65492 107936 65504
rect 107988 65492 107994 65544
rect 162210 65492 162216 65544
rect 162268 65532 162274 65544
rect 203058 65532 203064 65544
rect 162268 65504 203064 65532
rect 162268 65492 162274 65504
rect 203058 65492 203064 65504
rect 203116 65492 203122 65544
rect 69290 65424 69296 65476
rect 69348 65464 69354 65476
rect 155862 65464 155868 65476
rect 69348 65436 155868 65464
rect 69348 65424 69354 65436
rect 155862 65424 155868 65436
rect 155920 65424 155926 65476
rect 164142 65424 164148 65476
rect 164200 65464 164206 65476
rect 182634 65464 182640 65476
rect 164200 65436 182640 65464
rect 164200 65424 164206 65436
rect 182634 65424 182640 65436
rect 182692 65424 182698 65476
rect 68738 65356 68744 65408
rect 68796 65396 68802 65408
rect 109770 65396 109776 65408
rect 68796 65368 109776 65396
rect 68796 65356 68802 65368
rect 109770 65356 109776 65368
rect 109828 65356 109834 65408
rect 110874 65356 110880 65408
rect 110932 65396 110938 65408
rect 175826 65396 175832 65408
rect 110932 65368 175832 65396
rect 110932 65356 110938 65368
rect 175826 65356 175832 65368
rect 175884 65356 175890 65408
rect 73338 65288 73344 65340
rect 73396 65328 73402 65340
rect 106274 65328 106280 65340
rect 73396 65300 106280 65328
rect 73396 65288 73402 65300
rect 106274 65288 106280 65300
rect 106332 65288 106338 65340
rect 155862 65288 155868 65340
rect 155920 65328 155926 65340
rect 164878 65328 164884 65340
rect 155920 65300 164884 65328
rect 155920 65288 155926 65300
rect 164878 65288 164884 65300
rect 164936 65288 164942 65340
rect 90634 65220 90640 65272
rect 90692 65260 90698 65272
rect 125318 65260 125324 65272
rect 90692 65232 125324 65260
rect 90692 65220 90698 65232
rect 125318 65220 125324 65232
rect 125376 65220 125382 65272
rect 66162 64812 66168 64864
rect 66220 64852 66226 64864
rect 168282 64852 168288 64864
rect 66220 64824 168288 64852
rect 66220 64812 66226 64824
rect 168282 64812 168288 64824
rect 168340 64812 168346 64864
rect 66070 64744 66076 64796
rect 66128 64784 66134 64796
rect 167730 64784 167736 64796
rect 66128 64756 167736 64784
rect 66128 64744 66134 64756
rect 167730 64744 167736 64756
rect 167788 64744 167794 64796
rect 67542 64676 67548 64728
rect 67600 64716 67606 64728
rect 167454 64716 167460 64728
rect 67600 64688 167460 64716
rect 67600 64676 67606 64688
rect 167454 64676 167460 64688
rect 167512 64676 167518 64728
rect 69474 64608 69480 64660
rect 69532 64648 69538 64660
rect 168190 64648 168196 64660
rect 69532 64620 168196 64648
rect 69532 64608 69538 64620
rect 168190 64608 168196 64620
rect 168248 64608 168254 64660
rect 69750 64540 69756 64592
rect 69808 64580 69814 64592
rect 166994 64580 167000 64592
rect 69808 64552 167000 64580
rect 69808 64540 69814 64552
rect 166994 64540 167000 64552
rect 167052 64540 167058 64592
rect 69658 64472 69664 64524
rect 69716 64512 69722 64524
rect 168098 64512 168104 64524
rect 69716 64484 168104 64512
rect 69716 64472 69722 64484
rect 168098 64472 168104 64484
rect 168156 64472 168162 64524
rect 69842 64336 69848 64388
rect 69900 64376 69906 64388
rect 166074 64376 166080 64388
rect 69900 64348 166080 64376
rect 69900 64336 69906 64348
rect 166074 64336 166080 64348
rect 166132 64336 166138 64388
rect 168834 64336 168840 64388
rect 168892 64376 168898 64388
rect 249794 64376 249800 64388
rect 168892 64348 249800 64376
rect 168892 64336 168898 64348
rect 249794 64336 249800 64348
rect 249852 64336 249858 64388
rect 81710 64268 81716 64320
rect 81768 64308 81774 64320
rect 111058 64308 111064 64320
rect 81768 64280 111064 64308
rect 81768 64268 81774 64280
rect 111058 64268 111064 64280
rect 111116 64268 111122 64320
rect 168926 64268 168932 64320
rect 168984 64308 168990 64320
rect 270494 64308 270500 64320
rect 168984 64280 270500 64308
rect 168984 64268 168990 64280
rect 270494 64268 270500 64280
rect 270552 64268 270558 64320
rect 69382 64200 69388 64252
rect 69440 64240 69446 64252
rect 167638 64240 167644 64252
rect 69440 64212 167644 64240
rect 69440 64200 69446 64212
rect 167638 64200 167644 64212
rect 167696 64200 167702 64252
rect 169294 64200 169300 64252
rect 169352 64240 169358 64252
rect 285674 64240 285680 64252
rect 169352 64212 285680 64240
rect 169352 64200 169358 64212
rect 285674 64200 285680 64212
rect 285732 64200 285738 64252
rect 168098 64132 168104 64184
rect 168156 64172 168162 64184
rect 320174 64172 320180 64184
rect 168156 64144 320180 64172
rect 168156 64132 168162 64144
rect 320174 64132 320180 64144
rect 320232 64132 320238 64184
rect 110322 64064 110328 64116
rect 110380 64104 110386 64116
rect 196618 64104 196624 64116
rect 110380 64076 196624 64104
rect 110380 64064 110386 64076
rect 196618 64064 196624 64076
rect 196676 64064 196682 64116
rect 166074 63588 166080 63640
rect 166132 63628 166138 63640
rect 170398 63628 170404 63640
rect 166132 63600 170404 63628
rect 166132 63588 166138 63600
rect 170398 63588 170404 63600
rect 170456 63588 170462 63640
rect 167454 63520 167460 63572
rect 167512 63560 167518 63572
rect 169938 63560 169944 63572
rect 167512 63532 169944 63560
rect 167512 63520 167518 63532
rect 169938 63520 169944 63532
rect 169996 63520 170002 63572
rect 169570 62908 169576 62960
rect 169628 62948 169634 62960
rect 262214 62948 262220 62960
rect 169628 62920 262220 62948
rect 169628 62908 169634 62920
rect 262214 62908 262220 62920
rect 262272 62908 262278 62960
rect 166994 62840 167000 62892
rect 167052 62880 167058 62892
rect 288434 62880 288440 62892
rect 167052 62852 288440 62880
rect 167052 62840 167058 62852
rect 288434 62840 288440 62852
rect 288492 62840 288498 62892
rect 169018 62772 169024 62824
rect 169076 62812 169082 62824
rect 327074 62812 327080 62824
rect 169076 62784 327080 62812
rect 169076 62772 169082 62784
rect 327074 62772 327080 62784
rect 327132 62772 327138 62824
rect 169846 61480 169852 61532
rect 169904 61520 169910 61532
rect 242894 61520 242900 61532
rect 169904 61492 242900 61520
rect 169904 61480 169910 61492
rect 242894 61480 242900 61492
rect 242952 61480 242958 61532
rect 169386 61412 169392 61464
rect 169444 61452 169450 61464
rect 259546 61452 259552 61464
rect 169444 61424 259552 61452
rect 169444 61412 169450 61424
rect 259546 61412 259552 61424
rect 259604 61412 259610 61464
rect 167822 61344 167828 61396
rect 167880 61384 167886 61396
rect 307018 61384 307024 61396
rect 167880 61356 307024 61384
rect 167880 61344 167886 61356
rect 307018 61344 307024 61356
rect 307076 61344 307082 61396
rect 203610 60664 203616 60716
rect 203668 60704 203674 60716
rect 580166 60704 580172 60716
rect 203668 60676 580172 60704
rect 203668 60664 203674 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 168190 60052 168196 60104
rect 168248 60092 168254 60104
rect 248414 60092 248420 60104
rect 168248 60064 248420 60092
rect 168248 60052 168254 60064
rect 248414 60052 248420 60064
rect 248472 60052 248478 60104
rect 169938 59984 169944 60036
rect 169996 60024 170002 60036
rect 291194 60024 291200 60036
rect 169996 59996 291200 60024
rect 169996 59984 170002 59996
rect 291194 59984 291200 59996
rect 291252 59984 291258 60036
rect 196618 58624 196624 58676
rect 196676 58664 196682 58676
rect 284294 58664 284300 58676
rect 196676 58636 284300 58664
rect 196676 58624 196682 58636
rect 284294 58624 284300 58636
rect 284352 58624 284358 58676
rect 169202 57196 169208 57248
rect 169260 57236 169266 57248
rect 273254 57236 273260 57248
rect 169260 57208 273260 57236
rect 169260 57196 169266 57208
rect 273254 57196 273260 57208
rect 273312 57196 273318 57248
rect 170490 55904 170496 55956
rect 170548 55944 170554 55956
rect 264238 55944 264244 55956
rect 170548 55916 264244 55944
rect 170548 55904 170554 55916
rect 264238 55904 264244 55916
rect 264296 55904 264302 55956
rect 169110 55836 169116 55888
rect 169168 55876 169174 55888
rect 298094 55876 298100 55888
rect 169168 55848 298100 55876
rect 169168 55836 169174 55848
rect 298094 55836 298100 55848
rect 298152 55836 298158 55888
rect 194410 51688 194416 51740
rect 194468 51728 194474 51740
rect 333974 51728 333980 51740
rect 194468 51700 333980 51728
rect 194468 51688 194474 51700
rect 333974 51688 333980 51700
rect 334032 51688 334038 51740
rect 168282 50328 168288 50380
rect 168340 50368 168346 50380
rect 251266 50368 251272 50380
rect 168340 50340 251272 50368
rect 168340 50328 168346 50340
rect 251266 50328 251272 50340
rect 251324 50328 251330 50380
rect 178034 49036 178040 49088
rect 178092 49076 178098 49088
rect 245654 49076 245660 49088
rect 178092 49048 245660 49076
rect 178092 49036 178098 49048
rect 245654 49036 245660 49048
rect 245712 49036 245718 49088
rect 169478 48968 169484 49020
rect 169536 49008 169542 49020
rect 281534 49008 281540 49020
rect 169536 48980 281540 49008
rect 169536 48968 169542 48980
rect 281534 48968 281540 48980
rect 281592 48968 281598 49020
rect 171870 47540 171876 47592
rect 171928 47580 171934 47592
rect 345014 47580 345020 47592
rect 171928 47552 345020 47580
rect 171928 47540 171934 47552
rect 345014 47540 345020 47552
rect 345072 47540 345078 47592
rect 164878 46860 164884 46912
rect 164936 46900 164942 46912
rect 580166 46900 580172 46912
rect 164936 46872 580172 46900
rect 164936 46860 164942 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 186958 46180 186964 46232
rect 187016 46220 187022 46232
rect 247034 46220 247040 46232
rect 187016 46192 247040 46220
rect 187016 46180 187022 46192
rect 247034 46180 247040 46192
rect 247092 46180 247098 46232
rect 2774 45500 2780 45552
rect 2832 45540 2838 45552
rect 4798 45540 4804 45552
rect 2832 45512 4804 45540
rect 2832 45500 2838 45512
rect 4798 45500 4804 45512
rect 4856 45500 4862 45552
rect 170398 44820 170404 44872
rect 170456 44860 170462 44872
rect 292666 44860 292672 44872
rect 170456 44832 292672 44860
rect 170456 44820 170462 44832
rect 292666 44820 292672 44832
rect 292724 44820 292730 44872
rect 167730 42032 167736 42084
rect 167788 42072 167794 42084
rect 310514 42072 310520 42084
rect 167788 42044 310520 42072
rect 167788 42032 167794 42044
rect 310514 42032 310520 42044
rect 310572 42032 310578 42084
rect 167638 39312 167644 39364
rect 167696 39352 167702 39364
rect 269114 39352 269120 39364
rect 167696 39324 269120 39352
rect 167696 39312 167702 39324
rect 269114 39312 269120 39324
rect 269172 39312 269178 39364
rect 194502 37884 194508 37936
rect 194560 37924 194566 37936
rect 287054 37924 287060 37936
rect 194560 37896 287060 37924
rect 194560 37884 194566 37896
rect 287054 37884 287060 37896
rect 287112 37884 287118 37936
rect 171778 33736 171784 33788
rect 171836 33776 171842 33788
rect 311158 33776 311164 33788
rect 171836 33748 311164 33776
rect 171836 33736 171842 33748
rect 311158 33736 311164 33748
rect 311216 33736 311222 33788
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 65518 33096 65524 33108
rect 2924 33068 65524 33096
rect 2924 33056 2930 33068
rect 65518 33056 65524 33068
rect 65576 33056 65582 33108
rect 191098 33056 191104 33108
rect 191156 33096 191162 33108
rect 580166 33096 580172 33108
rect 191156 33068 580172 33096
rect 191156 33056 191162 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 190362 31016 190368 31068
rect 190420 31056 190426 31068
rect 322934 31056 322940 31068
rect 190420 31028 322940 31056
rect 190420 31016 190426 31028
rect 322934 31016 322940 31028
rect 322992 31016 322998 31068
rect 167270 28228 167276 28280
rect 167328 28268 167334 28280
rect 280154 28268 280160 28280
rect 167328 28240 280160 28268
rect 167328 28228 167334 28240
rect 280154 28228 280160 28240
rect 280212 28228 280218 28280
rect 169754 24080 169760 24132
rect 169812 24120 169818 24132
rect 263594 24120 263600 24132
rect 169812 24092 263600 24120
rect 169812 24080 169818 24092
rect 263594 24080 263600 24092
rect 263652 24080 263658 24132
rect 220078 22720 220084 22772
rect 220136 22760 220142 22772
rect 316126 22760 316132 22772
rect 220136 22732 316132 22760
rect 220136 22720 220142 22732
rect 316126 22720 316132 22732
rect 316184 22720 316190 22772
rect 198642 21360 198648 21412
rect 198700 21400 198706 21412
rect 266354 21400 266360 21412
rect 198700 21372 266360 21400
rect 198700 21360 198706 21372
rect 266354 21360 266360 21372
rect 266412 21360 266418 21412
rect 3510 20612 3516 20664
rect 3568 20652 3574 20664
rect 106366 20652 106372 20664
rect 3568 20624 106372 20652
rect 3568 20612 3574 20624
rect 106366 20612 106372 20624
rect 106424 20612 106430 20664
rect 188338 18572 188344 18624
rect 188396 18612 188402 18624
rect 278774 18612 278780 18624
rect 188396 18584 278780 18612
rect 188396 18572 188402 18584
rect 278774 18572 278780 18584
rect 278832 18572 278838 18624
rect 209038 17212 209044 17264
rect 209096 17252 209102 17264
rect 276014 17252 276020 17264
rect 209096 17224 276020 17252
rect 209096 17212 209102 17224
rect 276014 17212 276020 17224
rect 276072 17212 276078 17264
rect 169662 15852 169668 15904
rect 169720 15892 169726 15904
rect 301498 15892 301504 15904
rect 169720 15864 301504 15892
rect 169720 15852 169726 15864
rect 301498 15852 301504 15864
rect 301556 15852 301562 15904
rect 173158 14424 173164 14476
rect 173216 14464 173222 14476
rect 258258 14464 258264 14476
rect 173216 14436 258264 14464
rect 173216 14424 173222 14436
rect 258258 14424 258264 14436
rect 258316 14424 258322 14476
rect 167914 13064 167920 13116
rect 167972 13104 167978 13116
rect 284386 13104 284392 13116
rect 167972 13076 284392 13104
rect 167972 13064 167978 13076
rect 284386 13064 284392 13076
rect 284444 13064 284450 13116
rect 175918 11704 175924 11756
rect 175976 11744 175982 11756
rect 240134 11744 240140 11756
rect 175976 11716 240140 11744
rect 175976 11704 175982 11716
rect 240134 11704 240140 11716
rect 240192 11704 240198 11756
rect 259454 11704 259460 11756
rect 259512 11744 259518 11756
rect 260650 11744 260656 11756
rect 259512 11716 260656 11744
rect 259512 11704 259518 11716
rect 260650 11704 260656 11716
rect 260708 11704 260714 11756
rect 185578 7624 185584 7676
rect 185636 7664 185642 7676
rect 242986 7664 242992 7676
rect 185636 7636 242992 7664
rect 185636 7624 185642 7636
rect 242986 7624 242992 7636
rect 243044 7624 243050 7676
rect 206278 7556 206284 7608
rect 206336 7596 206342 7608
rect 277118 7596 277124 7608
rect 206336 7568 277124 7596
rect 206336 7556 206342 7568
rect 277118 7556 277124 7568
rect 277176 7556 277182 7608
rect 182818 6808 182824 6860
rect 182876 6848 182882 6860
rect 580166 6848 580172 6860
rect 182876 6820 580172 6848
rect 182876 6808 182882 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 187602 4972 187608 5024
rect 187660 5012 187666 5024
rect 274818 5012 274824 5024
rect 187660 4984 274824 5012
rect 187660 4972 187666 4984
rect 274818 4972 274824 4984
rect 274876 4972 274882 5024
rect 180058 4904 180064 4956
rect 180116 4944 180122 4956
rect 322106 4944 322112 4956
rect 180116 4916 322112 4944
rect 180116 4904 180122 4916
rect 322106 4904 322112 4916
rect 322164 4904 322170 4956
rect 181438 4836 181444 4888
rect 181496 4876 181502 4888
rect 324406 4876 324412 4888
rect 181496 4848 324412 4876
rect 181496 4836 181502 4848
rect 324406 4836 324412 4848
rect 324464 4836 324470 4888
rect 4154 4768 4160 4820
rect 4212 4808 4218 4820
rect 107654 4808 107660 4820
rect 4212 4780 107660 4808
rect 4212 4768 4218 4780
rect 107654 4768 107660 4780
rect 107712 4768 107718 4820
rect 174538 4768 174544 4820
rect 174596 4808 174602 4820
rect 343358 4808 343364 4820
rect 174596 4780 343364 4808
rect 174596 4768 174602 4780
rect 343358 4768 343364 4780
rect 343416 4768 343422 4820
rect 238726 3828 248414 3856
rect 235258 3680 235264 3732
rect 235316 3720 235322 3732
rect 238726 3720 238754 3828
rect 245194 3788 245200 3800
rect 235316 3692 238754 3720
rect 241992 3760 245200 3788
rect 235316 3680 235322 3692
rect 177390 3612 177396 3664
rect 177448 3652 177454 3664
rect 241992 3652 242020 3760
rect 245194 3748 245200 3760
rect 245252 3748 245258 3800
rect 248386 3720 248414 3828
rect 267734 3720 267740 3732
rect 248386 3692 267740 3720
rect 267734 3680 267740 3692
rect 267792 3680 267798 3732
rect 177448 3624 242020 3652
rect 177448 3612 177454 3624
rect 242894 3612 242900 3664
rect 242952 3652 242958 3664
rect 244090 3652 244096 3664
rect 242952 3624 244096 3652
rect 242952 3612 242958 3624
rect 244090 3612 244096 3624
rect 244148 3612 244154 3664
rect 251174 3612 251180 3664
rect 251232 3652 251238 3664
rect 252370 3652 252376 3664
rect 251232 3624 252376 3652
rect 251232 3612 251238 3624
rect 252370 3612 252376 3624
rect 252428 3612 252434 3664
rect 284294 3612 284300 3664
rect 284352 3652 284358 3664
rect 285030 3652 285036 3664
rect 284352 3624 285036 3652
rect 284352 3612 284358 3624
rect 285030 3612 285036 3624
rect 285088 3612 285094 3664
rect 299566 3612 299572 3664
rect 299624 3652 299630 3664
rect 300762 3652 300768 3664
rect 299624 3624 300768 3652
rect 299624 3612 299630 3624
rect 300762 3612 300768 3624
rect 300820 3612 300826 3664
rect 311158 3612 311164 3664
rect 311216 3652 311222 3664
rect 312630 3652 312636 3664
rect 311216 3624 312636 3652
rect 311216 3612 311222 3624
rect 312630 3612 312636 3624
rect 312688 3612 312694 3664
rect 203518 3544 203524 3596
rect 203576 3584 203582 3596
rect 319714 3584 319720 3596
rect 203576 3556 319720 3584
rect 203576 3544 203582 3556
rect 319714 3544 319720 3556
rect 319772 3544 319778 3596
rect 324314 3544 324320 3596
rect 324372 3584 324378 3596
rect 325602 3584 325608 3596
rect 324372 3556 325608 3584
rect 324372 3544 324378 3556
rect 325602 3544 325608 3556
rect 325660 3544 325666 3596
rect 332686 3544 332692 3596
rect 332744 3584 332750 3596
rect 333882 3584 333888 3596
rect 332744 3556 333888 3584
rect 332744 3544 332750 3556
rect 333882 3544 333888 3556
rect 333940 3544 333946 3596
rect 344554 3584 344560 3596
rect 335326 3556 344560 3584
rect 184198 3476 184204 3528
rect 184256 3516 184262 3528
rect 335326 3516 335354 3556
rect 344554 3544 344560 3556
rect 344612 3544 344618 3596
rect 184256 3488 335354 3516
rect 184256 3476 184262 3488
rect 340966 3476 340972 3528
rect 341024 3516 341030 3528
rect 342162 3516 342168 3528
rect 341024 3488 342168 3516
rect 341024 3476 341030 3488
rect 342162 3476 342168 3488
rect 342220 3476 342226 3528
rect 349154 3476 349160 3528
rect 349212 3516 349218 3528
rect 350442 3516 350448 3528
rect 349212 3488 350448 3516
rect 349212 3476 349218 3488
rect 350442 3476 350448 3488
rect 350500 3476 350506 3528
rect 69106 3408 69112 3460
rect 69164 3448 69170 3460
rect 136450 3448 136456 3460
rect 69164 3420 136456 3448
rect 69164 3408 69170 3420
rect 136450 3408 136456 3420
rect 136508 3408 136514 3460
rect 177298 3408 177304 3460
rect 177356 3448 177362 3460
rect 177356 3420 341012 3448
rect 177356 3408 177362 3420
rect 340984 3392 341012 3420
rect 307018 3340 307024 3392
rect 307076 3380 307082 3392
rect 309042 3380 309048 3392
rect 307076 3352 309048 3380
rect 307076 3340 307082 3352
rect 309042 3340 309048 3352
rect 309100 3340 309106 3392
rect 316034 3340 316040 3392
rect 316092 3380 316098 3392
rect 317322 3380 317328 3392
rect 316092 3352 317328 3380
rect 316092 3340 316098 3352
rect 317322 3340 317328 3352
rect 317380 3340 317386 3392
rect 340966 3340 340972 3392
rect 341024 3340 341030 3392
rect 264238 3136 264244 3188
rect 264296 3176 264302 3188
rect 265342 3176 265348 3188
rect 264296 3148 265348 3176
rect 264296 3136 264302 3148
rect 265342 3136 265348 3148
rect 265400 3136 265406 3188
rect 566 2796 572 2848
rect 624 2836 630 2848
rect 4154 2836 4160 2848
rect 624 2808 4160 2836
rect 624 2796 630 2808
rect 4154 2796 4160 2808
rect 4212 2796 4218 2848
<< via1 >>
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 188344 700476 188396 700528
rect 267648 700476 267700 700528
rect 40500 700408 40552 700460
rect 78680 700408 78732 700460
rect 89168 700408 89220 700460
rect 122840 700408 122892 700460
rect 184204 700408 184256 700460
rect 364984 700408 365036 700460
rect 73068 700340 73120 700392
rect 137836 700340 137888 700392
rect 182824 700340 182876 700392
rect 429844 700340 429896 700392
rect 8116 700272 8168 700324
rect 94504 700272 94556 700324
rect 105452 700272 105504 700324
rect 120724 700272 120776 700324
rect 186964 700272 187016 700324
rect 527180 700272 527232 700324
rect 24308 699660 24360 699712
rect 25504 699660 25556 699712
rect 66168 699660 66220 699712
rect 72976 699660 73028 699712
rect 396724 699660 396776 699712
rect 397460 699660 397512 699712
rect 3424 683136 3476 683188
rect 75920 683136 75972 683188
rect 233884 683136 233936 683188
rect 579620 683136 579672 683188
rect 3516 670692 3568 670744
rect 55864 670692 55916 670744
rect 192484 670692 192536 670744
rect 580172 670692 580224 670744
rect 3424 656888 3476 656940
rect 95884 656888 95936 656940
rect 249064 643084 249116 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 54484 632068 54536 632120
rect 239404 630640 239456 630692
rect 579988 630640 580040 630692
rect 3148 618264 3200 618316
rect 106280 618264 106332 618316
rect 235264 616836 235316 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 62764 605820 62816 605872
rect 242164 590656 242216 590708
rect 580172 590656 580224 590708
rect 3332 579640 3384 579692
rect 65524 579640 65576 579692
rect 169668 576852 169720 576904
rect 580172 576852 580224 576904
rect 3424 565836 3476 565888
rect 11704 565836 11756 565888
rect 233976 563048 234028 563100
rect 580172 563048 580224 563100
rect 3424 553392 3476 553444
rect 121460 553392 121512 553444
rect 278044 536800 278096 536852
rect 579896 536800 579948 536852
rect 3424 527144 3476 527196
rect 120816 527144 120868 527196
rect 3424 514768 3476 514820
rect 107660 514768 107712 514820
rect 173164 510620 173216 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 99380 500964 99432 501016
rect 169576 484372 169628 484424
rect 580172 484372 580224 484424
rect 2780 474784 2832 474836
rect 4804 474784 4856 474836
rect 289084 470568 289136 470620
rect 580172 470568 580224 470620
rect 3240 462340 3292 462392
rect 18604 462340 18656 462392
rect 203524 456764 203576 456816
rect 580172 456764 580224 456816
rect 3148 448536 3200 448588
rect 61384 448536 61436 448588
rect 3424 422288 3476 422340
rect 119344 422288 119396 422340
rect 169852 418140 169904 418192
rect 580172 418140 580224 418192
rect 180064 404336 180116 404388
rect 580172 404336 580224 404388
rect 3516 397468 3568 397520
rect 10324 397468 10376 397520
rect 238024 378156 238076 378208
rect 580172 378156 580224 378208
rect 244924 364352 244976 364404
rect 579804 364352 579856 364404
rect 234068 351908 234120 351960
rect 580172 351908 580224 351960
rect 3332 345040 3384 345092
rect 71780 345040 71832 345092
rect 195244 324300 195296 324352
rect 579620 324300 579672 324352
rect 3332 318792 3384 318844
rect 15844 318792 15896 318844
rect 169944 311856 169996 311908
rect 580172 311856 580224 311908
rect 169024 298120 169076 298172
rect 580172 298120 580224 298172
rect 3332 292544 3384 292596
rect 58624 292544 58676 292596
rect 3424 266364 3476 266416
rect 7564 266364 7616 266416
rect 123668 265616 123720 265668
rect 201500 265616 201552 265668
rect 3608 260108 3660 260160
rect 120172 260108 120224 260160
rect 3332 258680 3384 258732
rect 120356 258680 120408 258732
rect 228364 258068 228416 258120
rect 579988 258068 580040 258120
rect 25504 257320 25556 257372
rect 121920 257320 121972 257372
rect 167736 257320 167788 257372
rect 542360 257320 542412 257372
rect 10324 255960 10376 256012
rect 121736 255960 121788 256012
rect 170036 255960 170088 256012
rect 234620 255960 234672 256012
rect 65892 254736 65944 254788
rect 170036 254736 170088 254788
rect 104164 254668 104216 254720
rect 155224 254668 155276 254720
rect 91284 254600 91336 254652
rect 68744 254532 68796 254584
rect 126336 254532 126388 254584
rect 142896 254532 142948 254584
rect 194600 254532 194652 254584
rect 91928 254464 91980 254516
rect 151084 254464 151136 254516
rect 195980 254464 196032 254516
rect 67548 254396 67600 254448
rect 153200 254396 153252 254448
rect 153844 254396 153896 254448
rect 69296 254328 69348 254380
rect 167276 254328 167328 254380
rect 69020 254260 69072 254312
rect 167184 254260 167236 254312
rect 69388 254192 69440 254244
rect 167644 254192 167696 254244
rect 67456 254124 67508 254176
rect 167736 254124 167788 254176
rect 73896 254056 73948 254108
rect 173992 254056 174044 254108
rect 77760 253988 77812 254040
rect 179420 253988 179472 254040
rect 3148 253920 3200 253972
rect 10324 253920 10376 253972
rect 114468 253920 114520 253972
rect 126980 253920 127032 253972
rect 155224 253920 155276 253972
rect 211160 253920 211212 253972
rect 80980 253512 81032 253564
rect 183652 253512 183704 253564
rect 68468 253444 68520 253496
rect 124864 253444 124916 253496
rect 99012 253376 99064 253428
rect 204904 253376 204956 253428
rect 93216 253240 93268 253292
rect 126244 253240 126296 253292
rect 126888 253240 126940 253292
rect 85488 253172 85540 253224
rect 133328 253172 133380 253224
rect 68744 253104 68796 253156
rect 120908 253104 120960 253156
rect 93860 253036 93912 253088
rect 148324 253036 148376 253088
rect 198740 253036 198792 253088
rect 68284 252968 68336 253020
rect 124036 252968 124088 253020
rect 126888 252968 126940 253020
rect 181444 252968 181496 253020
rect 90640 252900 90692 252952
rect 164148 252900 164200 252952
rect 194692 252900 194744 252952
rect 111892 252832 111944 252884
rect 142804 252832 142856 252884
rect 219440 252832 219492 252884
rect 89352 252764 89404 252816
rect 165528 252764 165580 252816
rect 193220 252764 193272 252816
rect 69480 252696 69532 252748
rect 167828 252696 167880 252748
rect 112536 252628 112588 252680
rect 121000 252628 121052 252680
rect 103520 252560 103572 252612
rect 119988 252560 120040 252612
rect 109960 252220 110012 252272
rect 118056 252220 118108 252272
rect 105452 252152 105504 252204
rect 118792 252152 118844 252204
rect 80336 252084 80388 252136
rect 112168 252084 112220 252136
rect 113180 252084 113232 252136
rect 124220 252084 124272 252136
rect 69204 252016 69256 252068
rect 71780 252016 71832 252068
rect 72608 252016 72660 252068
rect 121368 252016 121420 252068
rect 102232 251948 102284 252000
rect 157984 251948 158036 252000
rect 71320 251880 71372 251932
rect 122104 251880 122156 251932
rect 75828 251812 75880 251864
rect 130384 251812 130436 251864
rect 108028 251744 108080 251796
rect 124312 251744 124364 251796
rect 101588 251676 101640 251728
rect 125140 251676 125192 251728
rect 66076 251608 66128 251660
rect 75920 251608 75972 251660
rect 76472 251608 76524 251660
rect 95148 251608 95200 251660
rect 97080 251608 97132 251660
rect 127808 251608 127860 251660
rect 62028 251540 62080 251592
rect 85488 251540 85540 251592
rect 86776 251540 86828 251592
rect 124128 251540 124180 251592
rect 63408 251472 63460 251524
rect 74540 251472 74592 251524
rect 122196 251472 122248 251524
rect 117044 251404 117096 251456
rect 126704 251404 126756 251456
rect 61752 251336 61804 251388
rect 80980 251336 81032 251388
rect 110604 251336 110656 251388
rect 121276 251336 121328 251388
rect 157984 251336 158036 251388
rect 177304 251336 177356 251388
rect 97724 251268 97776 251320
rect 103428 251268 103480 251320
rect 118332 251268 118384 251320
rect 144184 251268 144236 251320
rect 211068 251268 211120 251320
rect 61936 251200 61988 251252
rect 75828 251200 75880 251252
rect 100300 251200 100352 251252
rect 117228 251200 117280 251252
rect 118976 251200 119028 251252
rect 126612 251200 126664 251252
rect 131120 251200 131172 251252
rect 131856 251200 131908 251252
rect 222844 251200 222896 251252
rect 107660 251132 107712 251184
rect 108672 251132 108724 251184
rect 203064 251132 203116 251184
rect 203524 251132 203576 251184
rect 211068 251132 211120 251184
rect 227720 251132 227772 251184
rect 228364 251132 228416 251184
rect 117964 250724 118016 250776
rect 125048 250724 125100 250776
rect 68192 250656 68244 250708
rect 123852 250656 123904 250708
rect 108672 250588 108724 250640
rect 134524 250588 134576 250640
rect 95884 250520 95936 250572
rect 117228 250520 117280 250572
rect 129740 250520 129792 250572
rect 130476 250452 130528 250504
rect 82912 250384 82964 250436
rect 121092 250384 121144 250436
rect 68008 250316 68060 250368
rect 123944 250316 123996 250368
rect 68652 250248 68704 250300
rect 124956 250248 125008 250300
rect 68836 250180 68888 250232
rect 117964 250180 118016 250232
rect 67916 250044 67968 250096
rect 127716 250112 127768 250164
rect 87420 250044 87472 250096
rect 146944 250112 146996 250164
rect 190460 250112 190512 250164
rect 152464 250044 152516 250096
rect 203064 250044 203116 250096
rect 63316 249976 63368 250028
rect 82912 249976 82964 250028
rect 99656 249976 99708 250028
rect 121184 249976 121236 250028
rect 129740 249976 129792 250028
rect 130568 249976 130620 250028
rect 205732 249976 205784 250028
rect 68376 249908 68428 249960
rect 123484 249908 123536 249960
rect 130476 249908 130528 249960
rect 201500 249908 201552 249960
rect 106740 249840 106792 249892
rect 140044 249840 140096 249892
rect 210424 249840 210476 249892
rect 64788 249772 64840 249824
rect 78680 249772 78732 249824
rect 79232 249772 79284 249824
rect 119804 249772 119856 249824
rect 134524 249772 134576 249824
rect 215944 249772 215996 249824
rect 118700 249704 118752 249756
rect 187700 249704 187752 249756
rect 188344 249704 188396 249756
rect 119160 249636 119212 249688
rect 119436 249636 119488 249688
rect 115480 249500 115532 249552
rect 119160 249500 119212 249552
rect 118056 249432 118108 249484
rect 118792 249432 118844 249484
rect 67088 249092 67140 249144
rect 67548 249092 67600 249144
rect 119712 249092 119764 249144
rect 121552 249092 121604 249144
rect 156604 249092 156656 249144
rect 159364 249024 159416 249076
rect 119712 248956 119764 249008
rect 119988 248956 120040 249008
rect 156604 248616 156656 248668
rect 212540 248616 212592 248668
rect 68744 248548 68796 248600
rect 126428 248548 126480 248600
rect 159364 248548 159416 248600
rect 218152 248548 218204 248600
rect 119160 248480 119212 248532
rect 69848 248412 69900 248464
rect 126520 248412 126572 248464
rect 162124 248412 162176 248464
rect 223580 248412 223632 248464
rect 121460 248344 121512 248396
rect 121828 248344 121880 248396
rect 119252 247732 119304 247784
rect 127624 247732 127676 247784
rect 10324 247664 10376 247716
rect 67640 247664 67692 247716
rect 119896 247664 119948 247716
rect 172612 247664 172664 247716
rect 127624 247188 127676 247240
rect 200120 247188 200172 247240
rect 133788 247120 133840 247172
rect 213368 247120 213420 247172
rect 121460 247052 121512 247104
rect 230296 247052 230348 247104
rect 121368 246440 121420 246492
rect 173900 246440 173952 246492
rect 122196 246372 122248 246424
rect 175464 246372 175516 246424
rect 122012 246304 122064 246356
rect 122380 246304 122432 246356
rect 229468 246304 229520 246356
rect 122656 245692 122708 245744
rect 129004 245692 129056 245744
rect 121460 245624 121512 245676
rect 122012 245624 122064 245676
rect 230204 245624 230256 245676
rect 121276 244944 121328 244996
rect 137284 244944 137336 244996
rect 15844 244876 15896 244928
rect 64512 244876 64564 244928
rect 122104 244876 122156 244928
rect 171140 244876 171192 244928
rect 137284 244468 137336 244520
rect 218060 244468 218112 244520
rect 121460 244400 121512 244452
rect 230940 244400 230992 244452
rect 121644 244332 121696 244384
rect 231308 244332 231360 244384
rect 64512 244264 64564 244316
rect 67640 244264 67692 244316
rect 205640 244264 205692 244316
rect 580172 244264 580224 244316
rect 68192 243584 68244 243636
rect 68836 243584 68888 243636
rect 68376 243516 68428 243568
rect 68652 243516 68704 243568
rect 66996 243448 67048 243500
rect 69480 243448 69532 243500
rect 122288 242972 122340 243024
rect 230112 242972 230164 243024
rect 121552 242904 121604 242956
rect 122104 242904 122156 242956
rect 231952 242904 232004 242956
rect 168288 242156 168340 242208
rect 205640 242156 205692 242208
rect 121552 241544 121604 241596
rect 230020 241544 230072 241596
rect 121460 241476 121512 241528
rect 231032 241476 231084 241528
rect 67088 240932 67140 240984
rect 68376 240932 68428 240984
rect 125140 240728 125192 240780
rect 159456 240728 159508 240780
rect 177304 240728 177356 240780
rect 208952 240728 209004 240780
rect 3056 240116 3108 240168
rect 66904 240116 66956 240168
rect 159456 240116 159508 240168
rect 207664 240116 207716 240168
rect 121828 239436 121880 239488
rect 147588 239436 147640 239488
rect 124128 239368 124180 239420
rect 158076 239368 158128 239420
rect 168932 239368 168984 239420
rect 282920 239368 282972 239420
rect 158076 238824 158128 238876
rect 190644 238824 190696 238876
rect 147588 238756 147640 238808
rect 231216 238756 231268 238808
rect 127808 237532 127860 237584
rect 131948 237532 132000 237584
rect 202880 237532 202932 237584
rect 121828 237464 121880 237516
rect 230756 237464 230808 237516
rect 121368 237328 121420 237380
rect 231124 237396 231176 237448
rect 130384 236784 130436 236836
rect 177120 236784 177172 236836
rect 186136 236784 186188 236836
rect 195244 236784 195296 236836
rect 129004 236716 129056 236768
rect 232688 236716 232740 236768
rect 169116 236648 169168 236700
rect 580356 236648 580408 236700
rect 122748 235968 122800 236020
rect 230572 235968 230624 236020
rect 126704 234744 126756 234796
rect 133236 234744 133288 234796
rect 226708 234744 226760 234796
rect 122288 234676 122340 234728
rect 229560 234676 229612 234728
rect 122472 234608 122524 234660
rect 230480 234608 230532 234660
rect 190460 233928 190512 233980
rect 191012 233928 191064 233980
rect 194600 233928 194652 233980
rect 195428 233928 195480 233980
rect 218060 233928 218112 233980
rect 218612 233928 218664 233980
rect 68468 233860 68520 233912
rect 68744 233860 68796 233912
rect 126612 233860 126664 233912
rect 229284 233860 229336 233912
rect 122472 233248 122524 233300
rect 230388 233248 230440 233300
rect 121276 233180 121328 233232
rect 122012 233180 122064 233232
rect 121092 233112 121144 233164
rect 186136 233180 186188 233232
rect 215944 233180 215996 233232
rect 217048 233180 217100 233232
rect 119344 233044 119396 233096
rect 171232 233112 171284 233164
rect 180064 233112 180116 233164
rect 210424 233112 210476 233164
rect 214472 233112 214524 233164
rect 213368 233044 213420 233096
rect 331220 233180 331272 233232
rect 222844 233112 222896 233164
rect 226064 233112 226116 233164
rect 121184 232772 121236 232824
rect 134616 232772 134668 232824
rect 119712 232704 119764 232756
rect 138664 232704 138716 232756
rect 121000 232636 121052 232688
rect 166816 232636 166868 232688
rect 66628 232568 66680 232620
rect 68744 232568 68796 232620
rect 133328 232568 133380 232620
rect 189356 232636 189408 232688
rect 181444 232568 181496 232620
rect 119804 232500 119856 232552
rect 181628 232500 181680 232552
rect 198372 232500 198424 232552
rect 226064 232500 226116 232552
rect 412640 232500 412692 232552
rect 166908 232092 166960 232144
rect 215760 232092 215812 232144
rect 140780 232024 140832 232076
rect 141424 232024 141476 232076
rect 192576 232024 192628 232076
rect 204904 232024 204956 232076
rect 234620 232024 234672 232076
rect 166816 231956 166868 232008
rect 221556 231956 221608 232008
rect 223488 231956 223540 232008
rect 233240 231956 233292 232008
rect 134616 231888 134668 231940
rect 206100 231888 206152 231940
rect 138664 231820 138716 231872
rect 210608 231820 210660 231872
rect 222200 231820 222252 231872
rect 234712 231820 234764 231872
rect 173992 231208 174044 231260
rect 175188 231208 175240 231260
rect 126520 231072 126572 231124
rect 150440 231072 150492 231124
rect 168196 231072 168248 231124
rect 579988 231072 580040 231124
rect 121736 230868 121788 230920
rect 122288 230868 122340 230920
rect 229100 230868 229152 230920
rect 121460 230800 121512 230852
rect 230664 230800 230716 230852
rect 169300 230732 169352 230784
rect 179420 230732 179472 230784
rect 169208 230664 169260 230716
rect 182456 230664 182508 230716
rect 150440 230596 150492 230648
rect 65800 230460 65852 230512
rect 67640 230460 67692 230512
rect 170036 230596 170088 230648
rect 183560 230596 183612 230648
rect 184848 230596 184900 230648
rect 198372 230596 198424 230648
rect 235356 230596 235408 230648
rect 169392 230528 169444 230580
rect 173992 230528 174044 230580
rect 65892 230392 65944 230444
rect 67732 230392 67784 230444
rect 169484 230460 169536 230512
rect 171140 230460 171192 230512
rect 170680 230392 170732 230444
rect 173164 230392 173216 230444
rect 229928 230392 229980 230444
rect 231952 230392 232004 230444
rect 163504 229848 163556 229900
rect 232320 229848 232372 229900
rect 120908 229780 120960 229832
rect 167000 229780 167052 229832
rect 166264 229712 166316 229764
rect 231952 229712 232004 229764
rect 166356 229644 166408 229696
rect 232136 229644 232188 229696
rect 166448 229576 166500 229628
rect 232228 229576 232280 229628
rect 166724 229508 166776 229560
rect 232504 229508 232556 229560
rect 166540 229440 166592 229492
rect 232412 229440 232464 229492
rect 165436 229372 165488 229424
rect 232596 229372 232648 229424
rect 162400 229304 162452 229356
rect 232044 229304 232096 229356
rect 144276 229168 144328 229220
rect 231860 229168 231912 229220
rect 121460 229100 121512 229152
rect 229284 229100 229336 229152
rect 229376 229100 229428 229152
rect 230848 229100 230900 229152
rect 125048 229032 125100 229084
rect 167092 229032 167144 229084
rect 231032 229032 231084 229084
rect 231400 229032 231452 229084
rect 233976 229032 234028 229084
rect 164884 226312 164936 226364
rect 167552 226312 167604 226364
rect 229652 226312 229704 226364
rect 548616 226312 548668 226364
rect 63500 225564 63552 225616
rect 64604 225564 64656 225616
rect 67824 225564 67876 225616
rect 122472 225564 122524 225616
rect 165436 225564 165488 225616
rect 66904 225292 66956 225344
rect 68744 225292 68796 225344
rect 15844 224952 15896 225004
rect 63500 224952 63552 225004
rect 119896 224952 119948 225004
rect 121552 224952 121604 225004
rect 139400 224952 139452 225004
rect 167092 224952 167144 225004
rect 121460 224884 121512 224936
rect 166724 224884 166776 224936
rect 124036 224816 124088 224868
rect 167092 224816 167144 224868
rect 230940 223524 230992 223576
rect 558920 223524 558972 223576
rect 125048 222164 125100 222216
rect 167092 222164 167144 222216
rect 121460 222028 121512 222080
rect 123668 222028 123720 222080
rect 124956 221416 125008 221468
rect 167460 221416 167512 221468
rect 65616 220804 65668 220856
rect 68008 220804 68060 220856
rect 120448 220736 120500 220788
rect 166540 220736 166592 220788
rect 67456 219444 67508 219496
rect 68928 219444 68980 219496
rect 119528 219376 119580 219428
rect 163504 219376 163556 219428
rect 235356 219376 235408 219428
rect 580172 219376 580224 219428
rect 153844 219308 153896 219360
rect 167092 219308 167144 219360
rect 119160 218424 119212 218476
rect 119528 218424 119580 218476
rect 120724 218084 120776 218136
rect 121552 218084 121604 218136
rect 65892 218016 65944 218068
rect 68192 218016 68244 218068
rect 121000 218016 121052 218068
rect 121460 218016 121512 218068
rect 119436 217948 119488 218000
rect 167092 217948 167144 218000
rect 232688 217948 232740 218000
rect 233884 217948 233936 218000
rect 122012 217268 122064 217320
rect 166448 217268 166500 217320
rect 66812 216656 66864 216708
rect 68376 216656 68428 216708
rect 121460 215976 121512 216028
rect 148416 215976 148468 216028
rect 123760 215908 123812 215960
rect 162860 215908 162912 215960
rect 167092 215908 167144 215960
rect 64420 215296 64472 215348
rect 67640 215296 67692 215348
rect 3332 215228 3384 215280
rect 15844 215228 15896 215280
rect 123944 214616 123996 214668
rect 144920 214616 144972 214668
rect 145932 214616 145984 214668
rect 3792 214548 3844 214600
rect 67640 214548 67692 214600
rect 123852 214548 123904 214600
rect 154580 214548 154632 214600
rect 155684 214548 155736 214600
rect 120816 214004 120868 214056
rect 121552 214004 121604 214056
rect 155684 214004 155736 214056
rect 167184 214004 167236 214056
rect 121460 213936 121512 213988
rect 142988 213936 143040 213988
rect 145932 213936 145984 213988
rect 167092 213936 167144 213988
rect 121736 213868 121788 213920
rect 144276 213868 144328 213920
rect 119988 212848 120040 212900
rect 122104 212848 122156 212900
rect 121920 212508 121972 212560
rect 156788 212508 156840 212560
rect 121184 212440 121236 212492
rect 122472 212440 122524 212492
rect 121460 211760 121512 211812
rect 122012 211760 122064 211812
rect 166356 211760 166408 211812
rect 121460 211624 121512 211676
rect 121920 211624 121972 211676
rect 162216 211488 162268 211540
rect 167092 211488 167144 211540
rect 162308 210808 162360 210860
rect 167092 210808 167144 210860
rect 123576 209720 123628 209772
rect 168196 209720 168248 209772
rect 230388 209720 230440 209772
rect 234068 209720 234120 209772
rect 229836 208360 229888 208412
rect 230388 208360 230440 208412
rect 124864 207612 124916 207664
rect 158720 207612 158772 207664
rect 158720 207000 158772 207052
rect 167092 207000 167144 207052
rect 548616 206932 548668 206984
rect 579988 206932 580040 206984
rect 137928 206388 137980 206440
rect 167092 206388 167144 206440
rect 121552 206320 121604 206372
rect 122104 206320 122156 206372
rect 162400 206320 162452 206372
rect 123484 206252 123536 206304
rect 167092 206252 167144 206304
rect 67364 205640 67416 205692
rect 68376 205640 68428 205692
rect 121092 205640 121144 205692
rect 122288 205640 122340 205692
rect 232688 205640 232740 205692
rect 548524 205640 548576 205692
rect 11704 205572 11756 205624
rect 67824 205572 67876 205624
rect 68008 204892 68060 204944
rect 69388 204892 69440 204944
rect 122564 204892 122616 204944
rect 166264 204892 166316 204944
rect 65708 204280 65760 204332
rect 68100 204280 68152 204332
rect 119804 204280 119856 204332
rect 121460 204280 121512 204332
rect 233148 204280 233200 204332
rect 580264 204280 580316 204332
rect 232688 204212 232740 204264
rect 278044 204212 278096 204264
rect 126428 203532 126480 203584
rect 167276 203532 167328 203584
rect 122564 202852 122616 202904
rect 164976 202852 165028 202904
rect 232688 202784 232740 202836
rect 289084 202784 289136 202836
rect 126336 202104 126388 202156
rect 167460 202104 167512 202156
rect 3424 201492 3476 201544
rect 63500 201492 63552 201544
rect 66720 201492 66772 201544
rect 67640 201492 67692 201544
rect 121828 201492 121880 201544
rect 124404 201492 124456 201544
rect 127716 201424 127768 201476
rect 167092 201424 167144 201476
rect 167276 201152 167328 201204
rect 167276 200948 167328 201000
rect 233332 200744 233384 200796
rect 477500 200744 477552 200796
rect 69388 200336 69440 200388
rect 72608 200336 72660 200388
rect 69848 200268 69900 200320
rect 71274 200268 71326 200320
rect 73252 200268 73304 200320
rect 74540 200268 74592 200320
rect 67180 200132 67232 200184
rect 69756 200132 69808 200184
rect 4804 200064 4856 200116
rect 7564 199996 7616 200048
rect 69572 199996 69624 200048
rect 75184 200268 75236 200320
rect 76472 200268 76524 200320
rect 77116 200268 77168 200320
rect 77760 200268 77812 200320
rect 79048 200268 79100 200320
rect 79692 200268 79744 200320
rect 80980 200268 81032 200320
rect 81624 200268 81676 200320
rect 82912 200268 82964 200320
rect 83556 200268 83608 200320
rect 84200 200268 84252 200320
rect 85488 200268 85540 200320
rect 86132 200268 86184 200320
rect 87420 200268 87472 200320
rect 88064 200268 88116 200320
rect 89352 200268 89404 200320
rect 89996 200268 90048 200320
rect 90640 200268 90692 200320
rect 91928 200268 91980 200320
rect 92572 200268 92624 200320
rect 93860 200268 93912 200320
rect 94504 200268 94556 200320
rect 95792 200268 95844 200320
rect 96436 200268 96488 200320
rect 97724 200268 97776 200320
rect 98368 200268 98420 200320
rect 102830 200336 102882 200388
rect 99012 200268 99064 200320
rect 100300 200268 100352 200320
rect 100898 200268 100950 200320
rect 102232 200268 102284 200320
rect 104164 200268 104216 200320
rect 73160 199928 73212 199980
rect 73252 199928 73304 199980
rect 74540 199928 74592 199980
rect 75092 199928 75144 199980
rect 76472 199928 76524 199980
rect 77116 199928 77168 199980
rect 77760 199928 77812 199980
rect 79048 199928 79100 199980
rect 79692 199928 79744 199980
rect 80980 199928 81032 199980
rect 81624 199928 81676 199980
rect 82912 199928 82964 199980
rect 83556 199928 83608 199980
rect 84200 199928 84252 199980
rect 85488 199928 85540 199980
rect 86132 199928 86184 199980
rect 87420 199928 87472 199980
rect 87972 199928 88024 199980
rect 89352 199928 89404 199980
rect 89904 199928 89956 199980
rect 90640 199928 90692 199980
rect 91836 199928 91888 199980
rect 92480 199928 92532 199980
rect 93860 199928 93912 199980
rect 94412 199928 94464 199980
rect 95700 199928 95752 199980
rect 96436 199928 96488 199980
rect 97264 199928 97316 199980
rect 98276 199928 98328 199980
rect 98552 199928 98604 199980
rect 98920 199928 98972 199980
rect 100300 199928 100352 199980
rect 101312 199928 101364 199980
rect 111248 200336 111300 200388
rect 104808 200268 104860 200320
rect 105406 200268 105458 200320
rect 106740 200268 106792 200320
rect 107384 200268 107436 200320
rect 103428 199928 103480 199980
rect 104164 199928 104216 199980
rect 104256 199928 104308 199980
rect 104808 199928 104860 199980
rect 105360 199928 105412 199980
rect 64512 199860 64564 199912
rect 75184 199860 75236 199912
rect 84660 199860 84712 199912
rect 62764 199792 62816 199844
rect 61384 199724 61436 199776
rect 75276 199724 75328 199776
rect 84844 199792 84896 199844
rect 98644 199792 98696 199844
rect 108672 200268 108724 200320
rect 109316 200268 109368 200320
rect 110604 200268 110656 200320
rect 107476 199928 107528 199980
rect 108764 199928 108816 199980
rect 109316 199928 109368 199980
rect 111248 199928 111300 199980
rect 111156 199860 111208 199912
rect 113180 200336 113232 200388
rect 111892 200268 111944 200320
rect 113778 200268 113830 200320
rect 115112 200268 115164 200320
rect 115756 200268 115808 200320
rect 117044 200268 117096 200320
rect 117688 200268 117740 200320
rect 112536 199928 112588 199980
rect 113180 199928 113232 199980
rect 114468 199928 114520 199980
rect 115296 199928 115348 199980
rect 115848 199928 115900 199980
rect 116584 199928 116636 199980
rect 119160 200472 119212 200524
rect 122564 200132 122616 200184
rect 152556 200132 152608 200184
rect 119068 200064 119120 200116
rect 117320 199928 117372 199980
rect 117688 199928 117740 199980
rect 138020 199928 138072 199980
rect 98736 199724 98788 199776
rect 65524 199656 65576 199708
rect 74816 199656 74868 199708
rect 75000 199656 75052 199708
rect 107200 199792 107252 199844
rect 69572 199588 69624 199640
rect 74724 199588 74776 199640
rect 75276 199588 75328 199640
rect 112536 199724 112588 199776
rect 113824 199724 113876 199776
rect 125048 199724 125100 199776
rect 108120 199656 108172 199708
rect 120080 199656 120132 199708
rect 108672 199588 108724 199640
rect 120448 199588 120500 199640
rect 68744 199520 68796 199572
rect 157340 199520 157392 199572
rect 69020 199452 69072 199504
rect 167368 199452 167420 199504
rect 65616 199384 65668 199436
rect 168196 199384 168248 199436
rect 169024 199384 169076 199436
rect 67916 199316 67968 199368
rect 72700 199316 72752 199368
rect 73160 199316 73212 199368
rect 84752 199316 84804 199368
rect 84936 199316 84988 199368
rect 75184 199248 75236 199300
rect 82084 199248 82136 199300
rect 74724 199180 74776 199232
rect 84660 199180 84712 199232
rect 84752 199180 84804 199232
rect 98552 199248 98604 199300
rect 98736 199316 98788 199368
rect 113732 199316 113784 199368
rect 113824 199248 113876 199300
rect 98644 199180 98696 199232
rect 117688 199180 117740 199232
rect 65800 199112 65852 199164
rect 84844 199112 84896 199164
rect 117136 198908 117188 198960
rect 122380 198908 122432 198960
rect 117228 198840 117280 198892
rect 122012 198840 122064 198892
rect 117044 198772 117096 198824
rect 121644 198772 121696 198824
rect 68836 198704 68888 198756
rect 71044 198704 71096 198756
rect 118516 198704 118568 198756
rect 121552 198704 121604 198756
rect 68560 198636 68612 198688
rect 164884 198636 164936 198688
rect 18604 198568 18656 198620
rect 87420 198568 87472 198620
rect 91836 198568 91888 198620
rect 58624 198500 58676 198552
rect 104072 198500 104124 198552
rect 108764 198568 108816 198620
rect 110420 198568 110472 198620
rect 55864 198432 55916 198484
rect 97264 198432 97316 198484
rect 98920 198432 98972 198484
rect 106280 198432 106332 198484
rect 113824 198500 113876 198552
rect 117320 198500 117372 198552
rect 111800 198432 111852 198484
rect 66168 198364 66220 198416
rect 75092 198364 75144 198416
rect 81624 198364 81676 198416
rect 106924 198364 106976 198416
rect 107200 198364 107252 198416
rect 127072 198364 127124 198416
rect 101312 198296 101364 198348
rect 129740 198296 129792 198348
rect 104256 198228 104308 198280
rect 131120 198228 131172 198280
rect 65800 198160 65852 198212
rect 79048 198160 79100 198212
rect 95700 198160 95752 198212
rect 126336 198160 126388 198212
rect 63224 198092 63276 198144
rect 69388 198092 69440 198144
rect 107476 198092 107528 198144
rect 137284 198092 137336 198144
rect 157340 198092 157392 198144
rect 158168 198092 158220 198144
rect 167368 198092 167420 198144
rect 61844 198024 61896 198076
rect 79692 198024 79744 198076
rect 85488 198024 85540 198076
rect 111064 198024 111116 198076
rect 114468 198024 114520 198076
rect 170312 198024 170364 198076
rect 65892 197956 65944 198008
rect 168288 197956 168340 198008
rect 169760 197956 169812 198008
rect 86132 197888 86184 197940
rect 109040 197888 109092 197940
rect 77116 197820 77168 197872
rect 79324 197820 79376 197872
rect 89904 197820 89956 197872
rect 108396 197820 108448 197872
rect 104072 197752 104124 197804
rect 111156 197752 111208 197804
rect 104808 197684 104860 197736
rect 109132 197684 109184 197736
rect 104164 197616 104216 197668
rect 110512 197616 110564 197668
rect 137284 197616 137336 197668
rect 166356 197616 166408 197668
rect 131120 197548 131172 197600
rect 131764 197548 131816 197600
rect 166448 197548 166500 197600
rect 126336 197480 126388 197532
rect 166264 197480 166316 197532
rect 117964 197412 118016 197464
rect 119160 197412 119212 197464
rect 129740 197412 129792 197464
rect 130384 197412 130436 197464
rect 170404 197412 170456 197464
rect 92480 197344 92532 197396
rect 94596 197344 94648 197396
rect 118608 197344 118660 197396
rect 119620 197344 119672 197396
rect 127072 197344 127124 197396
rect 127716 197344 127768 197396
rect 170496 197344 170548 197396
rect 76472 196732 76524 196784
rect 86224 196732 86276 196784
rect 108764 196732 108816 196784
rect 119436 196732 119488 196784
rect 69112 196664 69164 196716
rect 128360 196664 128412 196716
rect 69480 196596 69532 196648
rect 70308 196596 70360 196648
rect 167368 196596 167420 196648
rect 118700 195984 118752 196036
rect 119712 195984 119764 196036
rect 169024 195984 169076 196036
rect 105360 195508 105412 195560
rect 113272 195508 113324 195560
rect 100300 195440 100352 195492
rect 110604 195440 110656 195492
rect 98276 195372 98328 195424
rect 113364 195372 113416 195424
rect 94412 195304 94464 195356
rect 115940 195304 115992 195356
rect 87972 195236 88024 195288
rect 114560 195236 114612 195288
rect 115664 194896 115716 194948
rect 121920 194896 121972 194948
rect 116584 194624 116636 194676
rect 166540 194624 166592 194676
rect 3424 194556 3476 194608
rect 117964 194556 118016 194608
rect 113088 193944 113140 193996
rect 118700 193944 118752 193996
rect 108488 193876 108540 193928
rect 120172 193876 120224 193928
rect 63500 193808 63552 193860
rect 111892 193808 111944 193860
rect 122104 193808 122156 193860
rect 115756 193672 115808 193724
rect 122748 193672 122800 193724
rect 68468 192448 68520 192500
rect 167368 192448 167420 192500
rect 233884 191836 233936 191888
rect 579712 191836 579764 191888
rect 66812 191088 66864 191140
rect 168104 191088 168156 191140
rect 233148 191088 233200 191140
rect 233424 191088 233476 191140
rect 578884 191088 578936 191140
rect 115848 190544 115900 190596
rect 113824 190476 113876 190528
rect 118056 190476 118108 190528
rect 162400 190476 162452 190528
rect 89352 189796 89404 189848
rect 123484 189796 123536 189848
rect 64420 189728 64472 189780
rect 155868 189728 155920 189780
rect 142988 189116 143040 189168
rect 144276 189116 144328 189168
rect 155868 189116 155920 189168
rect 167368 189116 167420 189168
rect 123484 189048 123536 189100
rect 164884 189048 164936 189100
rect 110236 188300 110288 188352
rect 122656 188300 122708 188352
rect 233148 188300 233200 188352
rect 233516 188300 233568 188352
rect 242164 188300 242216 188352
rect 72700 186940 72752 186992
rect 150532 186940 150584 186992
rect 233148 186940 233200 186992
rect 233608 186940 233660 186992
rect 249064 186940 249116 186992
rect 150532 186328 150584 186380
rect 151728 186328 151780 186380
rect 167368 186328 167420 186380
rect 69664 185580 69716 185632
rect 167368 185580 167420 185632
rect 68008 184832 68060 184884
rect 167368 184832 167420 184884
rect 82912 184152 82964 184204
rect 116676 184152 116728 184204
rect 116676 183540 116728 183592
rect 156880 183540 156932 183592
rect 72608 183472 72660 183524
rect 167368 183472 167420 183524
rect 110328 183404 110380 183456
rect 115296 183404 115348 183456
rect 117964 183404 118016 183456
rect 123852 183404 123904 183456
rect 90640 182792 90692 182844
rect 123484 182792 123536 182844
rect 123484 182180 123536 182232
rect 163504 182180 163556 182232
rect 77760 181432 77812 181484
rect 112444 181432 112496 181484
rect 112444 180820 112496 180872
rect 163596 180820 163648 180872
rect 71044 180072 71096 180124
rect 167460 180072 167512 180124
rect 97264 177352 97316 177404
rect 123208 177352 123260 177404
rect 68928 177284 68980 177336
rect 167460 177284 167512 177336
rect 123208 176672 123260 176724
rect 123668 176672 123720 176724
rect 166632 176672 166684 176724
rect 65708 175924 65760 175976
rect 69388 175924 69440 175976
rect 168104 175924 168156 175976
rect 233056 175176 233108 175228
rect 494060 175176 494112 175228
rect 111248 174496 111300 174548
rect 140780 174496 140832 174548
rect 140780 173884 140832 173936
rect 141516 173884 141568 173936
rect 168932 173884 168984 173936
rect 80980 173204 81032 173256
rect 114468 173204 114520 173256
rect 66720 173136 66772 173188
rect 168748 173136 168800 173188
rect 170312 173000 170364 173052
rect 170312 172796 170364 172848
rect 113916 172524 113968 172576
rect 114468 172524 114520 172576
rect 168748 172524 168800 172576
rect 68652 172456 68704 172508
rect 168104 172456 168156 172508
rect 112536 171912 112588 171964
rect 123760 171912 123812 171964
rect 111156 171844 111208 171896
rect 134708 171844 134760 171896
rect 70492 171776 70544 171828
rect 170404 171776 170456 171828
rect 231768 171776 231820 171828
rect 462320 171776 462372 171828
rect 134708 171164 134760 171216
rect 169852 171164 169904 171216
rect 123760 171096 123812 171148
rect 169576 171096 169628 171148
rect 231676 171028 231728 171080
rect 231952 171028 232004 171080
rect 170496 170824 170548 170876
rect 96436 170620 96488 170672
rect 125600 170620 125652 170672
rect 126888 170620 126940 170672
rect 170496 170620 170548 170672
rect 83556 170552 83608 170604
rect 115388 170552 115440 170604
rect 169852 170552 169904 170604
rect 109316 170484 109368 170536
rect 143448 170484 143500 170536
rect 75184 170416 75236 170468
rect 109224 170416 109276 170468
rect 69296 170348 69348 170400
rect 168104 170348 168156 170400
rect 169852 170348 169904 170400
rect 228824 170348 228876 170400
rect 231860 170348 231912 170400
rect 168656 170280 168708 170332
rect 173256 170280 173308 170332
rect 167920 170212 167972 170264
rect 171968 170212 172020 170264
rect 173900 170212 173952 170264
rect 175188 170212 175240 170264
rect 142988 169940 143040 169992
rect 143448 169940 143500 169992
rect 170404 170144 170456 170196
rect 126888 169872 126940 169924
rect 170036 170008 170088 170060
rect 176476 170212 176528 170264
rect 177764 170212 177816 170264
rect 178408 170212 178460 170264
rect 179696 170212 179748 170264
rect 180984 170212 181036 170264
rect 181628 170212 181680 170264
rect 182916 170212 182968 170264
rect 184204 170212 184256 170264
rect 185492 170212 185544 170264
rect 186136 170212 186188 170264
rect 187424 170212 187476 170264
rect 188712 170212 188764 170264
rect 189356 170212 189408 170264
rect 190644 170212 190696 170264
rect 191932 170212 191984 170264
rect 193220 170212 193272 170264
rect 193864 170212 193916 170264
rect 195152 170212 195204 170264
rect 196440 170212 196492 170264
rect 197084 170212 197136 170264
rect 198372 170212 198424 170264
rect 199660 170212 199712 170264
rect 200948 170212 201000 170264
rect 201592 170212 201644 170264
rect 202880 170212 202932 170264
rect 204168 170212 204220 170264
rect 204812 170212 204864 170264
rect 206100 170212 206152 170264
rect 207388 170212 207440 170264
rect 208676 170212 208728 170264
rect 209320 170212 209372 170264
rect 210608 170212 210660 170264
rect 211896 170212 211948 170264
rect 212540 170212 212592 170264
rect 213828 170212 213880 170264
rect 215116 170212 215168 170264
rect 216404 170212 216456 170264
rect 217048 170212 217100 170264
rect 218336 170212 218388 170264
rect 219624 170212 219676 170264
rect 220268 170212 220320 170264
rect 221556 170212 221608 170264
rect 222844 170212 222896 170264
rect 224132 170212 224184 170264
rect 224776 170212 224828 170264
rect 226064 170212 226116 170264
rect 227352 170212 227404 170264
rect 173900 169940 173952 169992
rect 175188 169940 175240 169992
rect 175280 169940 175332 169992
rect 177764 169940 177816 169992
rect 178408 169940 178460 169992
rect 179696 169940 179748 169992
rect 180984 169940 181036 169992
rect 181628 169940 181680 169992
rect 182916 169940 182968 169992
rect 184204 169940 184256 169992
rect 185492 169940 185544 169992
rect 186136 169940 186188 169992
rect 187424 169940 187476 169992
rect 188712 169940 188764 169992
rect 189356 169940 189408 169992
rect 189448 169940 189500 169992
rect 191932 169940 191984 169992
rect 193220 169940 193272 169992
rect 193864 169940 193916 169992
rect 195152 169940 195204 169992
rect 196440 169940 196492 169992
rect 196532 169940 196584 169992
rect 198372 169940 198424 169992
rect 199660 169940 199712 169992
rect 201408 169940 201460 169992
rect 201592 169940 201644 169992
rect 202880 169940 202932 169992
rect 204168 169940 204220 169992
rect 204812 169940 204864 169992
rect 206100 169940 206152 169992
rect 207388 169940 207440 169992
rect 208676 169940 208728 169992
rect 115388 169804 115440 169856
rect 170956 169872 171008 169924
rect 109224 169736 109276 169788
rect 109684 169736 109736 169788
rect 171048 169804 171100 169856
rect 168012 169736 168064 169788
rect 169668 169736 169720 169788
rect 166448 169668 166500 169720
rect 210608 169940 210660 169992
rect 211896 169940 211948 169992
rect 212540 169940 212592 169992
rect 213828 169940 213880 169992
rect 215116 169940 215168 169992
rect 216404 169940 216456 169992
rect 217048 169940 217100 169992
rect 218336 169940 218388 169992
rect 219624 169940 219676 169992
rect 220268 169940 220320 169992
rect 221556 169940 221608 169992
rect 222844 169940 222896 169992
rect 224776 169940 224828 169992
rect 226064 169940 226116 169992
rect 227352 169940 227404 169992
rect 115296 169600 115348 169652
rect 73252 169328 73304 169380
rect 108304 169532 108356 169584
rect 173900 169532 173952 169584
rect 175188 169532 175240 169584
rect 238024 169532 238076 169584
rect 166356 169464 166408 169516
rect 215116 169464 215168 169516
rect 118056 169396 118108 169448
rect 181168 169396 181220 169448
rect 198372 169396 198424 169448
rect 235264 169396 235316 169448
rect 170496 169328 170548 169380
rect 213828 169328 213880 169380
rect 79324 169260 79376 169312
rect 110696 169260 110748 169312
rect 170220 169260 170272 169312
rect 207388 169260 207440 169312
rect 94596 169192 94648 169244
rect 127808 169192 127860 169244
rect 196532 169192 196584 169244
rect 87604 169124 87656 169176
rect 122104 169124 122156 169176
rect 189448 169124 189500 169176
rect 84200 169056 84252 169108
rect 156696 169056 156748 169108
rect 169024 169056 169076 169108
rect 229284 169056 229336 169108
rect 103428 168988 103480 169040
rect 133328 168988 133380 169040
rect 208676 168988 208728 169040
rect 209688 168988 209740 169040
rect 580448 168988 580500 169040
rect 166264 168920 166316 168972
rect 201408 168920 201460 168972
rect 110696 168852 110748 168904
rect 111156 168852 111208 168904
rect 178408 168852 178460 168904
rect 184940 168852 184992 168904
rect 186136 168852 186188 168904
rect 396724 168852 396776 168904
rect 156696 168376 156748 168428
rect 187424 168376 187476 168428
rect 171048 168308 171100 168360
rect 175280 168308 175332 168360
rect 196440 168308 196492 168360
rect 203432 168308 203484 168360
rect 226064 168308 226116 168360
rect 347780 168308 347832 168360
rect 123852 168240 123904 168292
rect 228732 168240 228784 168292
rect 169576 168172 169628 168224
rect 220268 168172 220320 168224
rect 221556 168172 221608 168224
rect 299480 168172 299532 168224
rect 166632 168104 166684 168156
rect 202880 168104 202932 168156
rect 218336 168104 218388 168156
rect 239404 168104 239456 168156
rect 169852 168036 169904 168088
rect 219624 168036 219676 168088
rect 170404 167968 170456 168020
rect 217048 167968 217100 168020
rect 181168 167900 181220 167952
rect 227352 167900 227404 167952
rect 170036 167832 170088 167884
rect 201592 167832 201644 167884
rect 163504 167764 163556 167816
rect 195152 167764 195204 167816
rect 163964 167696 164016 167748
rect 168656 167696 168708 167748
rect 195244 167696 195296 167748
rect 233240 167696 233292 167748
rect 86224 167628 86276 167680
rect 111248 167628 111300 167680
rect 177764 167628 177816 167680
rect 195336 167628 195388 167680
rect 234712 167628 234764 167680
rect 164056 167560 164108 167612
rect 167920 167560 167972 167612
rect 189356 167560 189408 167612
rect 204352 167560 204404 167612
rect 162400 167492 162452 167544
rect 224776 167492 224828 167544
rect 163596 167424 163648 167476
rect 179696 167424 179748 167476
rect 193220 167424 193272 167476
rect 244924 167424 244976 167476
rect 156880 167356 156932 167408
rect 185492 167356 185544 167408
rect 182916 167288 182968 167340
rect 209688 167288 209740 167340
rect 548524 166948 548576 167000
rect 580172 166948 580224 167000
rect 226984 166404 227036 166456
rect 232228 166404 232280 166456
rect 215208 166336 215260 166388
rect 232504 166336 232556 166388
rect 202236 166268 202288 166320
rect 230020 166268 230072 166320
rect 108488 165520 108540 165572
rect 233424 165520 233476 165572
rect 108856 165452 108908 165504
rect 232412 165452 232464 165504
rect 108764 165384 108816 165436
rect 229560 165384 229612 165436
rect 121000 165316 121052 165368
rect 229376 165316 229428 165368
rect 111708 164908 111760 164960
rect 124404 165248 124456 165300
rect 231860 165248 231912 165300
rect 144276 165180 144328 165232
rect 144828 165180 144880 165232
rect 233516 165180 233568 165232
rect 148416 165112 148468 165164
rect 148968 165112 149020 165164
rect 232780 165112 232832 165164
rect 152556 165044 152608 165096
rect 153108 165044 153160 165096
rect 231952 165044 232004 165096
rect 164884 164976 164936 165028
rect 188712 164976 188764 165028
rect 209044 164976 209096 165028
rect 232688 164976 232740 165028
rect 166356 164908 166408 164960
rect 193864 164908 193916 164960
rect 202144 164908 202196 164960
rect 230940 164908 230992 164960
rect 119344 164840 119396 164892
rect 229468 164840 229520 164892
rect 166264 164772 166316 164824
rect 184204 164772 184256 164824
rect 163780 164704 163832 164756
rect 180984 164704 181036 164756
rect 163872 164636 163924 164688
rect 181628 164636 181680 164688
rect 224868 163548 224920 163600
rect 232044 163548 232096 163600
rect 164976 163480 165028 163532
rect 201500 163480 201552 163532
rect 231032 163480 231084 163532
rect 166724 162120 166776 162172
rect 191932 162120 191984 162172
rect 201408 162120 201460 162172
rect 580264 162120 580316 162172
rect 199936 160692 199988 160744
rect 230848 160692 230900 160744
rect 217968 159332 218020 159384
rect 229100 159332 229152 159384
rect 2964 149064 3016 149116
rect 106464 149064 106516 149116
rect 202328 142808 202380 142860
rect 231308 142808 231360 142860
rect 3516 137912 3568 137964
rect 61752 137912 61804 137964
rect 65524 137912 65576 137964
rect 220728 131724 220780 131776
rect 232596 131724 232648 131776
rect 119068 130228 119120 130280
rect 119620 130228 119672 130280
rect 201592 130364 201644 130416
rect 202236 130364 202288 130416
rect 122288 129004 122340 129056
rect 219440 129004 219492 129056
rect 220728 129004 220780 129056
rect 169668 127576 169720 127628
rect 580264 127576 580316 127628
rect 234620 126896 234672 126948
rect 580172 126896 580224 126948
rect 66996 126216 67048 126268
rect 169024 126216 169076 126268
rect 169668 126216 169720 126268
rect 183560 126216 183612 126268
rect 234620 126216 234672 126268
rect 147036 125468 147088 125520
rect 147588 125468 147640 125520
rect 162492 124992 162544 125044
rect 202236 124992 202288 125044
rect 162584 124924 162636 124976
rect 200488 124924 200540 124976
rect 111616 124856 111668 124908
rect 121460 124856 121512 124908
rect 147036 124856 147088 124908
rect 202052 124856 202104 124908
rect 119896 124788 119948 124840
rect 200028 124788 200080 124840
rect 121368 124720 121420 124772
rect 200396 124720 200448 124772
rect 121092 124652 121144 124704
rect 201776 124652 201828 124704
rect 119252 124584 119304 124636
rect 200304 124584 200356 124636
rect 121276 124516 121328 124568
rect 202880 124516 202932 124568
rect 119712 124448 119764 124500
rect 201684 124448 201736 124500
rect 115296 124380 115348 124432
rect 203156 124380 203208 124432
rect 108580 124312 108632 124364
rect 201868 124312 201920 124364
rect 108672 124244 108724 124296
rect 203064 124244 203116 124296
rect 174544 124176 174596 124228
rect 306380 124176 306432 124228
rect 109776 124108 109828 124160
rect 110236 124108 110288 124160
rect 119160 124108 119212 124160
rect 119528 124108 119580 124160
rect 120908 124108 120960 124160
rect 121184 124108 121236 124160
rect 164976 124108 165028 124160
rect 165528 124108 165580 124160
rect 182916 124108 182968 124160
rect 183560 124108 183612 124160
rect 202144 124108 202196 124160
rect 202420 124108 202472 124160
rect 208400 124108 208452 124160
rect 209044 124108 209096 124160
rect 167276 123700 167328 123752
rect 167828 123700 167880 123752
rect 165252 123632 165304 123684
rect 201960 123632 202012 123684
rect 229652 123632 229704 123684
rect 165160 123564 165212 123616
rect 202420 123564 202472 123616
rect 165068 123496 165120 123548
rect 202328 123496 202380 123548
rect 3424 123428 3476 123480
rect 95884 123428 95936 123480
rect 112536 123428 112588 123480
rect 112904 123428 112956 123480
rect 229100 123428 229152 123480
rect 229744 123428 229796 123480
rect 159548 123360 159600 123412
rect 205732 123360 205784 123412
rect 162400 123292 162452 123344
rect 208400 123292 208452 123344
rect 119528 123224 119580 123276
rect 200212 123224 200264 123276
rect 120908 123156 120960 123208
rect 204628 123156 204680 123208
rect 119436 123088 119488 123140
rect 164976 123088 165028 123140
rect 175832 123088 175884 123140
rect 259460 123088 259512 123140
rect 204536 123020 204588 123072
rect 115756 122952 115808 123004
rect 204720 122952 204772 123004
rect 112996 122884 113048 122936
rect 203248 122884 203300 122936
rect 109776 122816 109828 122868
rect 202972 122816 203024 122868
rect 170956 122612 171008 122664
rect 197728 122612 197780 122664
rect 179696 122544 179748 122596
rect 187700 122544 187752 122596
rect 155224 122476 155276 122528
rect 187424 122476 187476 122528
rect 88340 122408 88392 122460
rect 131948 122408 132000 122460
rect 181812 122408 181864 122460
rect 92204 122340 92256 122392
rect 130568 122340 130620 122392
rect 184756 122340 184808 122392
rect 99288 122272 99340 122324
rect 159364 122272 159416 122324
rect 93860 122204 93912 122256
rect 155224 122204 155276 122256
rect 163688 122272 163740 122324
rect 164148 122272 164200 122324
rect 173256 122272 173308 122324
rect 292580 122272 292632 122324
rect 191932 122204 191984 122256
rect 325700 122204 325752 122256
rect 91100 122136 91152 122188
rect 159456 122136 159508 122188
rect 185492 122136 185544 122188
rect 188068 122136 188120 122188
rect 198832 122136 198884 122188
rect 117136 122068 117188 122120
rect 226340 122068 226392 122120
rect 166816 122000 166868 122052
rect 193864 122000 193916 122052
rect 184756 121932 184808 121984
rect 200948 121932 201000 121984
rect 187424 121864 187476 121916
rect 203708 121864 203760 121916
rect 181812 121796 181864 121848
rect 200764 121796 200816 121848
rect 163688 121728 163740 121780
rect 175280 121728 175332 121780
rect 169760 121660 169812 121712
rect 186136 121728 186188 121780
rect 184848 121660 184900 121712
rect 190644 121660 190696 121712
rect 196440 121728 196492 121780
rect 206284 121728 206336 121780
rect 220084 121660 220136 121712
rect 226340 121660 226392 121712
rect 226984 121660 227036 121712
rect 104900 121592 104952 121644
rect 199016 121592 199068 121644
rect 199844 121592 199896 121644
rect 313280 121592 313332 121644
rect 186228 121524 186280 121576
rect 188068 121524 188120 121576
rect 116768 121456 116820 121508
rect 117136 121456 117188 121508
rect 169852 121456 169904 121508
rect 183560 121456 183612 121508
rect 186320 121456 186372 121508
rect 196440 121524 196492 121576
rect 193128 121456 193180 121508
rect 197084 121456 197136 121508
rect 102416 121388 102468 121440
rect 131120 121388 131172 121440
rect 143448 121388 143500 121440
rect 177120 121388 177172 121440
rect 103796 121320 103848 121372
rect 144184 121320 144236 121372
rect 148324 121320 148376 121372
rect 179696 121320 179748 121372
rect 95424 121252 95476 121304
rect 140044 121252 140096 121304
rect 190000 121252 190052 121304
rect 102140 121184 102192 121236
rect 162124 121184 162176 121236
rect 186320 121184 186372 121236
rect 83096 121116 83148 121168
rect 142896 121116 142948 121168
rect 143448 121116 143500 121168
rect 144184 121116 144236 121168
rect 198372 121116 198424 121168
rect 85580 121048 85632 121100
rect 148324 121048 148376 121100
rect 186228 121048 186280 121100
rect 94136 120980 94188 121032
rect 156604 120980 156656 121032
rect 158076 120980 158128 121032
rect 173256 120980 173308 121032
rect 80520 120912 80572 120964
rect 146944 120912 146996 120964
rect 174544 120912 174596 120964
rect 120724 120844 120776 120896
rect 227720 120844 227772 120896
rect 84200 120776 84252 120828
rect 151084 120776 151136 120828
rect 177764 120776 177816 120828
rect 86868 120708 86920 120760
rect 158076 120708 158128 120760
rect 187700 120776 187752 120828
rect 299480 120776 299532 120828
rect 305000 120708 305052 120760
rect 169760 120640 169812 120692
rect 184848 120640 184900 120692
rect 166172 120572 166224 120624
rect 195152 120572 195204 120624
rect 186780 120504 186832 120556
rect 203616 120504 203668 120556
rect 177120 120436 177172 120488
rect 203524 120436 203576 120488
rect 166080 120368 166132 120420
rect 195060 120368 195112 120420
rect 195796 120368 195848 120420
rect 227720 120368 227772 120420
rect 228732 120368 228784 120420
rect 168564 120300 168616 120352
rect 103612 119688 103664 119740
rect 133236 119960 133288 120012
rect 166448 120028 166500 120080
rect 169944 120232 169996 120284
rect 193864 120300 193916 120352
rect 252560 120300 252612 120352
rect 175280 120232 175332 120284
rect 176476 120232 176528 120284
rect 235264 120232 235316 120284
rect 182916 120164 182968 120216
rect 185492 120164 185544 120216
rect 295340 120164 295392 120216
rect 193220 120096 193272 120148
rect 580356 120096 580408 120148
rect 170956 120028 171008 120080
rect 135168 119892 135220 119944
rect 169760 119892 169812 119944
rect 169852 119892 169904 119944
rect 171968 119892 172020 119944
rect 199660 119892 199712 119944
rect 200580 119892 200632 119944
rect 86960 119620 87012 119672
rect 130476 119620 130528 119672
rect 166448 119824 166500 119876
rect 169116 119824 169168 119876
rect 171048 119824 171100 119876
rect 172428 119824 172480 119876
rect 197820 119824 197872 119876
rect 166632 119688 166684 119740
rect 166908 119688 166960 119740
rect 169668 119688 169720 119740
rect 89720 119552 89772 119604
rect 134616 119552 134668 119604
rect 135168 119552 135220 119604
rect 169852 119688 169904 119740
rect 79324 119484 79376 119536
rect 78496 119416 78548 119468
rect 78588 119348 78640 119400
rect 169116 119348 169168 119400
rect 198832 119824 198884 119876
rect 251180 119416 251232 119468
rect 271880 119348 271932 119400
rect 167276 119280 167328 119332
rect 169668 119280 169720 119332
rect 166448 118872 166500 118924
rect 200580 118940 200632 118992
rect 165344 118804 165396 118856
rect 200120 118804 200172 118856
rect 349160 118668 349212 118720
rect 64696 118600 64748 118652
rect 78496 118600 78548 118652
rect 138112 118600 138164 118652
rect 138664 118600 138716 118652
rect 164148 118600 164200 118652
rect 167184 118600 167236 118652
rect 167736 118600 167788 118652
rect 65984 118532 66036 118584
rect 77760 118532 77812 118584
rect 78588 118532 78640 118584
rect 157340 118532 157392 118584
rect 157984 118532 158036 118584
rect 169760 118532 169812 118584
rect 92480 118056 92532 118108
rect 138112 118056 138164 118108
rect 164792 118056 164844 118108
rect 165160 118056 165212 118108
rect 91560 117988 91612 118040
rect 157340 117988 157392 118040
rect 99840 117920 99892 117972
rect 166816 117920 166868 117972
rect 201960 117920 202012 117972
rect 202880 117920 202932 117972
rect 580264 117920 580316 117972
rect 80060 117444 80112 117496
rect 167092 117444 167144 117496
rect 75920 117376 75972 117428
rect 167000 117376 167052 117428
rect 65984 117308 66036 117360
rect 167920 117308 167972 117360
rect 63316 117240 63368 117292
rect 76472 117240 76524 117292
rect 77116 117240 77168 117292
rect 126244 117240 126296 117292
rect 126796 117240 126848 117292
rect 166540 117240 166592 117292
rect 64788 117172 64840 117224
rect 75920 117172 75972 117224
rect 137376 117172 137428 117224
rect 168656 117172 168708 117224
rect 98000 116696 98052 116748
rect 137376 116696 137428 116748
rect 84384 116628 84436 116680
rect 126796 116628 126848 116680
rect 82912 116560 82964 116612
rect 163688 116560 163740 116612
rect 202144 116560 202196 116612
rect 202972 116560 203024 116612
rect 282920 116560 282972 116612
rect 72608 116084 72660 116136
rect 169116 116084 169168 116136
rect 64420 116016 64472 116068
rect 167644 116016 167696 116068
rect 64696 115948 64748 116000
rect 167736 115948 167788 116000
rect 97724 115880 97776 115932
rect 99288 115880 99340 115932
rect 134616 115880 134668 115932
rect 165988 115880 166040 115932
rect 144920 115812 144972 115864
rect 145564 115812 145616 115864
rect 154580 115608 154632 115660
rect 155224 115608 155276 115660
rect 97080 115336 97132 115388
rect 134616 115336 134668 115388
rect 75552 115268 75604 115320
rect 80060 115268 80112 115320
rect 82268 115268 82320 115320
rect 164976 115268 165028 115320
rect 75828 115200 75880 115252
rect 166908 115200 166960 115252
rect 201960 115200 202012 115252
rect 203248 115200 203300 115252
rect 314660 115200 314712 115252
rect 64328 115064 64380 115116
rect 145564 115064 145616 115116
rect 69572 114996 69624 115048
rect 154580 114996 154632 115048
rect 73068 114928 73120 114980
rect 167000 114928 167052 114980
rect 71688 114860 71740 114912
rect 167184 114860 167236 114912
rect 66168 114792 66220 114844
rect 162860 114792 162912 114844
rect 163504 114792 163556 114844
rect 64236 114724 64288 114776
rect 162308 114724 162360 114776
rect 162676 114724 162728 114776
rect 70216 114656 70268 114708
rect 167092 114656 167144 114708
rect 65708 114588 65760 114640
rect 167828 114588 167880 114640
rect 64788 114520 64840 114572
rect 167552 114520 167604 114572
rect 60740 114452 60792 114504
rect 62028 114452 62080 114504
rect 79324 114452 79376 114504
rect 95884 114452 95936 114504
rect 96436 114452 96488 114504
rect 124312 114452 124364 114504
rect 166632 114452 166684 114504
rect 65524 114384 65576 114436
rect 75828 114384 75880 114436
rect 90640 114384 90692 114436
rect 92204 114384 92256 114436
rect 61936 114316 61988 114368
rect 71320 114316 71372 114368
rect 71688 114316 71740 114368
rect 74540 114316 74592 114368
rect 75920 114316 75972 114368
rect 67272 114248 67324 114300
rect 67548 114248 67600 114300
rect 100944 114248 100996 114300
rect 124220 114384 124272 114436
rect 166172 114384 166224 114436
rect 127624 114316 127676 114368
rect 168472 114316 168524 114368
rect 66076 114180 66128 114232
rect 71964 114180 72016 114232
rect 73068 114180 73120 114232
rect 101588 114180 101640 114232
rect 126980 114248 127032 114300
rect 166080 114248 166132 114300
rect 95148 114112 95200 114164
rect 133144 114180 133196 114232
rect 168380 114180 168432 114232
rect 86132 114044 86184 114096
rect 127624 114044 127676 114096
rect 99012 113976 99064 114028
rect 142804 113976 142856 114028
rect 143448 113976 143500 114028
rect 81624 113908 81676 113960
rect 140780 113908 140832 113960
rect 88708 113840 88760 113892
rect 152464 113840 152516 113892
rect 153016 113840 153068 113892
rect 3516 113772 3568 113824
rect 60740 113772 60792 113824
rect 64604 113772 64656 113824
rect 69388 113772 69440 113824
rect 89352 113772 89404 113824
rect 168564 113772 168616 113824
rect 200948 113772 201000 113824
rect 317420 113772 317472 113824
rect 79692 113636 79744 113688
rect 86868 113636 86920 113688
rect 70308 113568 70360 113620
rect 72332 113568 72384 113620
rect 67548 113500 67600 113552
rect 169116 113500 169168 113552
rect 72332 113432 72384 113484
rect 162308 113432 162360 113484
rect 69388 113364 69440 113416
rect 164976 113364 165028 113416
rect 68560 113296 68612 113348
rect 165528 113296 165580 113348
rect 64512 113228 64564 113280
rect 165344 113228 165396 113280
rect 166908 113160 166960 113212
rect 169300 113160 169352 113212
rect 200304 113228 200356 113280
rect 200212 113160 200264 113212
rect 202236 113092 202288 113144
rect 229928 113092 229980 113144
rect 200120 112820 200172 112872
rect 200212 112820 200264 112872
rect 69480 112480 69532 112532
rect 137928 112480 137980 112532
rect 71596 112412 71648 112464
rect 166908 112412 166960 112464
rect 67916 112344 67968 112396
rect 157984 112344 158036 112396
rect 68744 112276 68796 112328
rect 158720 112276 158772 112328
rect 69664 112208 69716 112260
rect 162216 112208 162268 112260
rect 68468 112140 68520 112192
rect 162124 112140 162176 112192
rect 67088 112072 67140 112124
rect 162768 112072 162820 112124
rect 65524 112004 65576 112056
rect 75184 112004 75236 112056
rect 75644 112004 75696 112056
rect 167000 112004 167052 112056
rect 70032 111936 70084 111988
rect 67088 111868 67140 111920
rect 67272 111868 67324 111920
rect 67824 111868 67876 111920
rect 68468 111868 68520 111920
rect 68928 111868 68980 111920
rect 70676 111868 70728 111920
rect 71596 111868 71648 111920
rect 169392 111936 169444 111988
rect 75460 111868 75512 111920
rect 101588 111868 101640 111920
rect 3424 111800 3476 111852
rect 100760 111800 100812 111852
rect 158720 111800 158772 111852
rect 159364 111800 159416 111852
rect 169392 111800 169444 111852
rect 169668 111800 169720 111852
rect 63408 111732 63460 111784
rect 68928 111732 68980 111784
rect 69296 111732 69348 111784
rect 70308 111732 70360 111784
rect 108948 111732 109000 111784
rect 111524 111732 111576 111784
rect 165252 111732 165304 111784
rect 69204 111664 69256 111716
rect 69848 111664 69900 111716
rect 75644 111664 75696 111716
rect 105728 111664 105780 111716
rect 119988 111664 120040 111716
rect 166448 111664 166500 111716
rect 108212 110508 108264 110560
rect 108580 110508 108632 110560
rect 70308 110440 70360 110492
rect 169484 110440 169536 110492
rect 108948 110372 109000 110424
rect 165160 110372 165212 110424
rect 202788 110372 202840 110424
rect 204720 110372 204772 110424
rect 108580 110304 108632 110356
rect 121276 110304 121328 110356
rect 150440 110304 150492 110356
rect 167000 110304 167052 110356
rect 201868 109760 201920 109812
rect 203156 109760 203208 109812
rect 267832 109760 267884 109812
rect 204720 109692 204772 109744
rect 299572 109692 299624 109744
rect 107660 108944 107712 108996
rect 109776 108944 109828 108996
rect 108028 108876 108080 108928
rect 116860 108944 116912 108996
rect 200304 108944 200356 108996
rect 200488 108944 200540 108996
rect 230572 108944 230624 108996
rect 231768 108944 231820 108996
rect 167552 108332 167604 108384
rect 167920 108332 167972 108384
rect 231768 108264 231820 108316
rect 336740 108264 336792 108316
rect 165528 107584 165580 107636
rect 167000 107584 167052 107636
rect 202788 107584 202840 107636
rect 205732 107584 205784 107636
rect 230480 107584 230532 107636
rect 231768 107584 231820 107636
rect 108948 107448 109000 107500
rect 164792 107448 164844 107500
rect 231768 106904 231820 106956
rect 347780 106904 347832 106956
rect 108948 106632 109000 106684
rect 112996 106632 113048 106684
rect 132500 106292 132552 106344
rect 167000 106292 167052 106344
rect 108948 106224 109000 106276
rect 165068 106224 165120 106276
rect 165344 106224 165396 106276
rect 167920 106224 167972 106276
rect 201868 105544 201920 105596
rect 230664 105544 230716 105596
rect 64512 104796 64564 104848
rect 67640 104796 67692 104848
rect 108028 104796 108080 104848
rect 119896 104796 119948 104848
rect 167460 104796 167512 104848
rect 169208 104796 169260 104848
rect 200764 104116 200816 104168
rect 289820 104116 289872 104168
rect 64788 103436 64840 103488
rect 67640 103436 67692 103488
rect 108948 103436 109000 103488
rect 147036 103436 147088 103488
rect 162032 103436 162084 103488
rect 167000 103436 167052 103488
rect 108212 103368 108264 103420
rect 121368 103368 121420 103420
rect 203708 102756 203760 102808
rect 255320 102756 255372 102808
rect 162768 102076 162820 102128
rect 167000 102076 167052 102128
rect 108948 102008 109000 102060
rect 115296 102008 115348 102060
rect 108580 101736 108632 101788
rect 108764 101736 108816 101788
rect 108764 101600 108816 101652
rect 115388 101600 115440 101652
rect 66076 100648 66128 100700
rect 67640 100648 67692 100700
rect 108948 100648 109000 100700
rect 162584 100648 162636 100700
rect 163504 100648 163556 100700
rect 167460 100648 167512 100700
rect 66168 100580 66220 100632
rect 68284 100580 68336 100632
rect 108764 100580 108816 100632
rect 159548 100580 159600 100632
rect 155224 100512 155276 100564
rect 167092 100512 167144 100564
rect 202788 100036 202840 100088
rect 208400 100036 208452 100088
rect 256700 100036 256752 100088
rect 201592 99968 201644 100020
rect 204628 99968 204680 100020
rect 307852 99968 307904 100020
rect 258724 99356 258776 99408
rect 580172 99356 580224 99408
rect 64328 99288 64380 99340
rect 67640 99288 67692 99340
rect 107660 99288 107712 99340
rect 162492 99288 162544 99340
rect 201592 99288 201644 99340
rect 219440 99288 219492 99340
rect 107752 98608 107804 98660
rect 119620 98608 119672 98660
rect 65984 97928 66036 97980
rect 67640 97928 67692 97980
rect 107660 97928 107712 97980
rect 121092 97928 121144 97980
rect 165528 97928 165580 97980
rect 166356 97928 166408 97980
rect 162216 97860 162268 97912
rect 167184 97860 167236 97912
rect 108396 96636 108448 96688
rect 165528 96636 165580 96688
rect 64236 96568 64288 96620
rect 67640 96568 67692 96620
rect 107844 96568 107896 96620
rect 119712 96568 119764 96620
rect 159364 96568 159416 96620
rect 168840 96568 168892 96620
rect 66628 96500 66680 96552
rect 69204 96500 69256 96552
rect 107660 96500 107712 96552
rect 119252 96500 119304 96552
rect 202144 95888 202196 95940
rect 203064 95888 203116 95940
rect 260840 95888 260892 95940
rect 107752 95208 107804 95260
rect 166448 95208 166500 95260
rect 201408 95208 201460 95260
rect 324320 95208 324372 95260
rect 107660 95140 107712 95192
rect 120080 95140 120132 95192
rect 120632 95140 120684 95192
rect 137928 95140 137980 95192
rect 167000 95140 167052 95192
rect 120080 94528 120132 94580
rect 166356 94528 166408 94580
rect 107660 94460 107712 94512
rect 119988 94460 120040 94512
rect 166540 94460 166592 94512
rect 202788 94460 202840 94512
rect 204536 94460 204588 94512
rect 296720 94460 296772 94512
rect 64696 93780 64748 93832
rect 67640 93780 67692 93832
rect 107752 93780 107804 93832
rect 162400 93780 162452 93832
rect 107660 93712 107712 93764
rect 120908 93712 120960 93764
rect 64420 92420 64472 92472
rect 67640 92420 67692 92472
rect 65708 92352 65760 92404
rect 68100 92352 68152 92404
rect 107752 91740 107804 91792
rect 122288 91740 122340 91792
rect 164976 90992 165028 91044
rect 167644 90992 167696 91044
rect 201776 90788 201828 90840
rect 204444 90788 204496 90840
rect 108028 90380 108080 90432
rect 120816 90380 120868 90432
rect 107660 90312 107712 90364
rect 119344 90312 119396 90364
rect 165068 90312 165120 90364
rect 204444 90312 204496 90364
rect 346400 90312 346452 90364
rect 201776 90040 201828 90092
rect 208400 90040 208452 90092
rect 107108 89700 107160 89752
rect 167000 89700 167052 89752
rect 157984 89632 158036 89684
rect 167184 89632 167236 89684
rect 202512 89632 202564 89684
rect 229100 89632 229152 89684
rect 230388 89632 230440 89684
rect 108580 88952 108632 89004
rect 166632 88952 166684 89004
rect 230388 88952 230440 89004
rect 329840 88952 329892 89004
rect 66904 88476 66956 88528
rect 68468 88476 68520 88528
rect 107292 88340 107344 88392
rect 167000 88340 167052 88392
rect 108948 88272 109000 88324
rect 119528 88272 119580 88324
rect 162308 88272 162360 88324
rect 167092 88272 167144 88324
rect 202512 88272 202564 88324
rect 226340 88272 226392 88324
rect 226800 88272 226852 88324
rect 226800 87592 226852 87644
rect 316040 87592 316092 87644
rect 3424 86980 3476 87032
rect 68100 86980 68152 87032
rect 67456 86912 67508 86964
rect 67916 86912 67968 86964
rect 108948 86912 109000 86964
rect 119436 86912 119488 86964
rect 164148 86912 164200 86964
rect 164884 86912 164936 86964
rect 202512 86912 202564 86964
rect 227812 86912 227864 86964
rect 227812 86232 227864 86284
rect 238760 86232 238812 86284
rect 200120 86096 200172 86148
rect 111064 85620 111116 85672
rect 164148 85620 164200 85672
rect 107200 85552 107252 85604
rect 167000 85552 167052 85604
rect 233884 85552 233936 85604
rect 580172 85552 580224 85604
rect 108212 85484 108264 85536
rect 144828 85484 144880 85536
rect 162124 85484 162176 85536
rect 167092 85484 167144 85536
rect 200120 85484 200172 85536
rect 3332 84804 3384 84856
rect 67640 84804 67692 84856
rect 67824 84804 67876 84856
rect 109224 84804 109276 84856
rect 122196 84804 122248 84856
rect 144828 84804 144880 84856
rect 164884 84804 164936 84856
rect 202696 84804 202748 84856
rect 203248 84804 203300 84856
rect 215208 84804 215260 84856
rect 277400 84804 277452 84856
rect 202696 84192 202748 84244
rect 203064 84192 203116 84244
rect 332600 84192 332652 84244
rect 108948 84124 109000 84176
rect 157248 84124 157300 84176
rect 157248 83512 157300 83564
rect 166816 83512 166868 83564
rect 155868 83444 155920 83496
rect 167000 83444 167052 83496
rect 203156 83444 203208 83496
rect 224868 83444 224920 83496
rect 331220 83444 331272 83496
rect 117228 82832 117280 82884
rect 162124 82832 162176 82884
rect 108948 82764 109000 82816
rect 67364 82356 67416 82408
rect 68468 82356 68520 82408
rect 108856 82084 108908 82136
rect 166908 82084 166960 82136
rect 107384 81404 107436 81456
rect 167000 81404 167052 81456
rect 108948 81336 109000 81388
rect 116768 81336 116820 81388
rect 108856 81268 108908 81320
rect 112536 81268 112588 81320
rect 151728 80656 151780 80708
rect 167000 80656 167052 80708
rect 107752 79976 107804 80028
rect 120724 79976 120776 80028
rect 166172 79296 166224 79348
rect 166724 79296 166776 79348
rect 202788 79296 202840 79348
rect 203340 79296 203392 79348
rect 217968 79296 218020 79348
rect 241520 79296 241572 79348
rect 108672 79228 108724 79280
rect 111892 79228 111944 79280
rect 118148 78752 118200 78804
rect 118516 78752 118568 78804
rect 164976 78752 165028 78804
rect 165160 78752 165212 78804
rect 167000 78752 167052 78804
rect 4804 78684 4856 78736
rect 65984 78684 66036 78736
rect 67640 78684 67692 78736
rect 106924 78684 106976 78736
rect 107936 78684 107988 78736
rect 166264 78684 166316 78736
rect 202788 78684 202840 78736
rect 204444 78684 204496 78736
rect 65432 78616 65484 78668
rect 66168 78616 66220 78668
rect 107752 78616 107804 78668
rect 118148 78616 118200 78668
rect 65340 78548 65392 78600
rect 66076 78548 66128 78600
rect 67640 78548 67692 78600
rect 66168 77596 66220 77648
rect 67640 77596 67692 77648
rect 107752 77188 107804 77240
rect 111616 77256 111668 77308
rect 162216 77256 162268 77308
rect 118148 76032 118200 76084
rect 118608 76032 118660 76084
rect 162400 76032 162452 76084
rect 107844 75964 107896 76016
rect 108120 75964 108172 76016
rect 162308 75964 162360 76016
rect 107752 75896 107804 75948
rect 162860 75896 162912 75948
rect 201316 75896 201368 75948
rect 253940 75896 253992 75948
rect 200948 75828 201000 75880
rect 222844 75828 222896 75880
rect 223488 75828 223540 75880
rect 107844 75216 107896 75268
rect 118148 75216 118200 75268
rect 107752 75148 107804 75200
rect 111708 75148 111760 75200
rect 166724 75148 166776 75200
rect 223488 75148 223540 75200
rect 302240 75148 302292 75200
rect 106188 74536 106240 74588
rect 167092 74536 167144 74588
rect 200488 74536 200540 74588
rect 339500 74536 339552 74588
rect 107752 74468 107804 74520
rect 153108 74468 153160 74520
rect 201960 74468 202012 74520
rect 221464 74468 221516 74520
rect 117964 73312 118016 73364
rect 164792 73312 164844 73364
rect 165528 73244 165580 73296
rect 167184 73244 167236 73296
rect 106096 73176 106148 73228
rect 167092 73176 167144 73228
rect 107752 73108 107804 73160
rect 117964 73108 118016 73160
rect 66720 72428 66772 72480
rect 68284 72428 68336 72480
rect 106096 71816 106148 71868
rect 106188 71816 106240 71868
rect 106096 71544 106148 71596
rect 107568 71748 107620 71800
rect 167092 71748 167144 71800
rect 108488 71680 108540 71732
rect 200304 71680 200356 71732
rect 201960 71680 202012 71732
rect 580172 71748 580224 71800
rect 108580 71612 108632 71664
rect 148968 71612 149020 71664
rect 200396 71612 200448 71664
rect 162860 71544 162912 71596
rect 201500 71544 201552 71596
rect 164884 71476 164936 71528
rect 201868 71476 201920 71528
rect 167460 71408 167512 71460
rect 168012 71408 168064 71460
rect 200488 71340 200540 71392
rect 201316 71340 201368 71392
rect 106004 70728 106056 70780
rect 198832 70660 198884 70712
rect 204812 70660 204864 70712
rect 198096 70592 198148 70644
rect 211896 71000 211948 71052
rect 3608 70320 3660 70372
rect 74540 70388 74592 70440
rect 75184 70388 75236 70440
rect 76472 70388 76524 70440
rect 70400 70252 70452 70304
rect 71274 70252 71326 70304
rect 71964 70252 72016 70304
rect 72608 70252 72660 70304
rect 73252 70252 73304 70304
rect 67548 70048 67600 70100
rect 70032 70048 70084 70100
rect 73896 70252 73948 70304
rect 71964 69912 72016 69964
rect 72608 69912 72660 69964
rect 73344 69912 73396 69964
rect 73988 69912 74040 69964
rect 65984 69844 66036 69896
rect 73712 69844 73764 69896
rect 82872 70320 82924 70372
rect 77116 70252 77168 70304
rect 77760 70252 77812 70304
rect 78404 70252 78456 70304
rect 79048 70252 79100 70304
rect 79692 70252 79744 70304
rect 80336 70252 80388 70304
rect 80980 70252 81032 70304
rect 81624 70252 81676 70304
rect 74540 69912 74592 69964
rect 75184 69912 75236 69964
rect 76564 69912 76616 69964
rect 77116 69912 77168 69964
rect 77760 69912 77812 69964
rect 78404 69912 78456 69964
rect 79048 69912 79100 69964
rect 79692 69912 79744 69964
rect 80428 69912 80480 69964
rect 81072 69912 81124 69964
rect 81716 69912 81768 69964
rect 83556 70252 83608 70304
rect 84200 70252 84252 70304
rect 100944 70320 100996 70372
rect 84860 70252 84912 70304
rect 85488 70252 85540 70304
rect 86132 70252 86184 70304
rect 86776 70252 86828 70304
rect 87420 70252 87472 70304
rect 88064 70252 88116 70304
rect 89352 70252 89404 70304
rect 89996 70252 90048 70304
rect 90640 70252 90692 70304
rect 91284 70252 91336 70304
rect 91928 70252 91980 70304
rect 92572 70252 92624 70304
rect 93216 70252 93268 70304
rect 93860 70252 93912 70304
rect 94520 70252 94572 70304
rect 95792 70252 95844 70304
rect 96436 70252 96488 70304
rect 97080 70252 97132 70304
rect 97724 70252 97776 70304
rect 98368 70252 98420 70304
rect 99012 70252 99064 70304
rect 99656 70252 99708 70304
rect 100300 70252 100352 70304
rect 82912 69912 82964 69964
rect 83648 69912 83700 69964
rect 84200 69912 84252 69964
rect 84936 69912 84988 69964
rect 85488 69912 85540 69964
rect 86132 69912 86184 69964
rect 86776 69912 86828 69964
rect 87420 69912 87472 69964
rect 88064 69912 88116 69964
rect 89352 69912 89404 69964
rect 102232 70252 102284 70304
rect 102876 70252 102928 70304
rect 166080 70388 166132 70440
rect 168012 70388 168064 70440
rect 103520 70252 103572 70304
rect 104180 70252 104232 70304
rect 104824 70252 104876 70304
rect 105468 70252 105520 70304
rect 106188 70252 106240 70304
rect 108028 70320 108080 70372
rect 200120 70320 200172 70372
rect 164792 70252 164844 70304
rect 204444 70252 204496 70304
rect 165160 70184 165212 70236
rect 165252 70184 165304 70236
rect 203248 70184 203300 70236
rect 110328 70116 110380 70168
rect 200396 70116 200448 70168
rect 108672 70048 108724 70100
rect 200028 70048 200080 70100
rect 115756 69980 115808 70032
rect 200488 69980 200540 70032
rect 94688 69912 94740 69964
rect 95792 69912 95844 69964
rect 96436 69912 96488 69964
rect 97080 69912 97132 69964
rect 97724 69912 97776 69964
rect 98368 69912 98420 69964
rect 99012 69912 99064 69964
rect 99656 69912 99708 69964
rect 100300 69912 100352 69964
rect 100944 69912 100996 69964
rect 102140 69912 102192 69964
rect 102232 69912 102284 69964
rect 102876 69912 102928 69964
rect 103152 69912 103204 69964
rect 103520 69912 103572 69964
rect 104624 69912 104676 69964
rect 165068 69912 165120 69964
rect 201776 69912 201828 69964
rect 84476 69844 84528 69896
rect 89904 69844 89956 69896
rect 89996 69844 90048 69896
rect 90640 69844 90692 69896
rect 91284 69844 91336 69896
rect 91928 69844 91980 69896
rect 92572 69844 92624 69896
rect 93216 69844 93268 69896
rect 93860 69844 93912 69896
rect 70308 69776 70360 69828
rect 75368 69776 75420 69828
rect 84016 69776 84068 69828
rect 68560 69708 68612 69760
rect 68376 69640 68428 69692
rect 75276 69708 75328 69760
rect 165528 69844 165580 69896
rect 166724 69844 166776 69896
rect 195244 69844 195296 69896
rect 107292 69776 107344 69828
rect 166540 69776 166592 69828
rect 201684 69844 201736 69896
rect 195428 69776 195480 69828
rect 202236 69776 202288 69828
rect 102140 69708 102192 69760
rect 106464 69708 106516 69760
rect 166448 69708 166500 69760
rect 201592 69708 201644 69760
rect 75276 69572 75328 69624
rect 75368 69572 75420 69624
rect 84016 69572 84068 69624
rect 166908 69640 166960 69692
rect 202144 69640 202196 69692
rect 202788 69640 202840 69692
rect 210608 69640 210660 69692
rect 73712 69504 73764 69556
rect 84476 69504 84528 69556
rect 89904 69572 89956 69624
rect 103152 69572 103204 69624
rect 166632 69572 166684 69624
rect 107108 69504 107160 69556
rect 202420 69504 202472 69556
rect 202696 69436 202748 69488
rect 206100 69436 206152 69488
rect 104624 69096 104676 69148
rect 113180 69096 113232 69148
rect 113548 69096 113600 69148
rect 106188 69028 106240 69080
rect 115756 69028 115808 69080
rect 166264 69028 166316 69080
rect 178040 69028 178092 69080
rect 179052 69028 179104 69080
rect 97724 68960 97776 69012
rect 104164 68960 104216 69012
rect 63224 68892 63276 68944
rect 71964 68892 72016 68944
rect 163964 68960 164016 69012
rect 171784 68960 171836 69012
rect 196624 68960 196676 69012
rect 202788 68960 202840 69012
rect 166264 68892 166316 68944
rect 184204 68892 184256 68944
rect 192576 68892 192628 68944
rect 202604 68892 202656 68944
rect 61844 68824 61896 68876
rect 77760 68824 77812 68876
rect 91928 68824 91980 68876
rect 95148 68824 95200 68876
rect 97080 68824 97132 68876
rect 109132 68824 109184 68876
rect 212540 68960 212592 69012
rect 213828 68960 213880 69012
rect 92572 68756 92624 68808
rect 106280 68756 106332 68808
rect 193220 68756 193272 68808
rect 197728 68756 197780 68808
rect 198648 68756 198700 68808
rect 65800 68688 65852 68740
rect 77116 68688 77168 68740
rect 163780 68688 163832 68740
rect 177396 68688 177448 68740
rect 76564 68620 76616 68672
rect 104072 68620 104124 68672
rect 104164 68620 104216 68672
rect 113272 68620 113324 68672
rect 198372 68688 198424 68740
rect 193864 68620 193916 68672
rect 194416 68620 194468 68672
rect 202696 68620 202748 68672
rect 93216 68552 93268 68604
rect 110604 68552 110656 68604
rect 81072 68484 81124 68536
rect 156696 68484 156748 68536
rect 181444 68484 181496 68536
rect 193220 68484 193272 68536
rect 194324 68484 194376 68536
rect 198832 68484 198884 68536
rect 86776 68416 86828 68468
rect 111800 68416 111852 68468
rect 187424 68416 187476 68468
rect 72608 68348 72660 68400
rect 108120 68348 108172 68400
rect 172980 68348 173032 68400
rect 213828 68348 213880 68400
rect 293960 68348 294012 68400
rect 96436 68280 96488 68332
rect 104164 68280 104216 68332
rect 104256 68280 104308 68332
rect 112444 68280 112496 68332
rect 175924 68280 175976 68332
rect 202604 68280 202656 68332
rect 204168 68280 204220 68332
rect 350540 68280 350592 68332
rect 86132 68212 86184 68264
rect 123576 68212 123628 68264
rect 186964 68212 187016 68264
rect 87420 68076 87472 68128
rect 127808 68076 127860 68128
rect 188344 68144 188396 68196
rect 70492 68008 70544 68060
rect 170496 68008 170548 68060
rect 170680 68008 170732 68060
rect 104164 67940 104216 67992
rect 110512 67940 110564 67992
rect 68836 67328 68888 67380
rect 106004 67532 106056 67584
rect 113088 67532 113140 67584
rect 200672 67532 200724 67584
rect 204444 67532 204496 67584
rect 233884 67532 233936 67584
rect 99656 67464 99708 67516
rect 110420 67464 110472 67516
rect 199384 67464 199436 67516
rect 215300 67464 215352 67516
rect 102876 67396 102928 67448
rect 2872 67260 2924 67312
rect 103980 67260 104032 67312
rect 80428 67192 80480 67244
rect 115204 67328 115256 67380
rect 115848 67328 115900 67380
rect 175832 67396 175884 67448
rect 258724 67396 258776 67448
rect 123760 67328 123812 67380
rect 200580 67328 200632 67380
rect 104164 67260 104216 67312
rect 106556 67260 106608 67312
rect 109040 67260 109092 67312
rect 182916 67260 182968 67312
rect 204444 67260 204496 67312
rect 82912 67124 82964 67176
rect 127624 67192 127676 67244
rect 199016 67192 199068 67244
rect 109040 67124 109092 67176
rect 109684 67124 109736 67176
rect 173900 67124 173952 67176
rect 187424 67124 187476 67176
rect 203432 67124 203484 67176
rect 95792 67056 95844 67108
rect 131764 67056 131816 67108
rect 196440 67056 196492 67108
rect 93860 66988 93912 67040
rect 130384 66988 130436 67040
rect 194508 66988 194560 67040
rect 99012 66920 99064 66972
rect 137284 66920 137336 66972
rect 199660 66920 199712 66972
rect 100300 66852 100352 66904
rect 142988 66852 143040 66904
rect 198740 66852 198792 66904
rect 215300 66852 215352 66904
rect 216404 66852 216456 66904
rect 349252 66852 349304 66904
rect 98368 66784 98420 66836
rect 127624 66784 127676 66836
rect 165436 66784 165488 66836
rect 185584 66784 185636 66836
rect 67824 66716 67876 66768
rect 107384 66716 107436 66768
rect 115848 66716 115900 66768
rect 180984 66716 181036 66768
rect 68928 66648 68980 66700
rect 106096 66648 106148 66700
rect 73988 66580 74040 66632
rect 109040 66580 109092 66632
rect 85488 66172 85540 66224
rect 108396 66172 108448 66224
rect 162124 66172 162176 66224
rect 208400 66172 208452 66224
rect 91284 66104 91336 66156
rect 123668 66104 123720 66156
rect 191932 66104 191984 66156
rect 83648 66036 83700 66088
rect 121460 66036 121512 66088
rect 125324 66036 125376 66088
rect 125508 66036 125560 66088
rect 191104 66036 191156 66088
rect 191288 66036 191340 66088
rect 94688 65968 94740 66020
rect 133328 65968 133380 66020
rect 133788 65968 133840 66020
rect 135168 65968 135220 66020
rect 200764 65968 200816 66020
rect 67916 65900 67968 65952
rect 107200 65900 107252 65952
rect 162308 65900 162360 65952
rect 203156 65900 203208 65952
rect 84936 65832 84988 65884
rect 123484 65832 123536 65884
rect 124128 65832 124180 65884
rect 126888 65832 126940 65884
rect 190000 65832 190052 65884
rect 75184 65764 75236 65816
rect 110880 65764 110932 65816
rect 111156 65764 111208 65816
rect 121460 65764 121512 65816
rect 122104 65764 122156 65816
rect 183560 65764 183612 65816
rect 89996 65696 90048 65748
rect 126336 65696 126388 65748
rect 126888 65696 126940 65748
rect 133788 65696 133840 65748
rect 195152 65696 195204 65748
rect 208400 65696 208452 65748
rect 209044 65696 209096 65748
rect 124128 65628 124180 65680
rect 184848 65628 184900 65680
rect 102232 65560 102284 65612
rect 134708 65560 134760 65612
rect 135168 65560 135220 65612
rect 162400 65560 162452 65612
rect 203340 65560 203392 65612
rect 79048 65492 79100 65544
rect 107936 65492 107988 65544
rect 162216 65492 162268 65544
rect 203064 65492 203116 65544
rect 69296 65424 69348 65476
rect 155868 65424 155920 65476
rect 164148 65424 164200 65476
rect 182640 65424 182692 65476
rect 68744 65356 68796 65408
rect 109776 65356 109828 65408
rect 110880 65356 110932 65408
rect 175832 65356 175884 65408
rect 73344 65288 73396 65340
rect 106280 65288 106332 65340
rect 155868 65288 155920 65340
rect 164884 65288 164936 65340
rect 90640 65220 90692 65272
rect 125324 65220 125376 65272
rect 66168 64812 66220 64864
rect 168288 64812 168340 64864
rect 66076 64744 66128 64796
rect 167736 64744 167788 64796
rect 67548 64676 67600 64728
rect 167460 64676 167512 64728
rect 69480 64608 69532 64660
rect 168196 64608 168248 64660
rect 69756 64540 69808 64592
rect 167000 64540 167052 64592
rect 69664 64472 69716 64524
rect 168104 64472 168156 64524
rect 69848 64336 69900 64388
rect 166080 64336 166132 64388
rect 168840 64336 168892 64388
rect 249800 64336 249852 64388
rect 81716 64268 81768 64320
rect 111064 64268 111116 64320
rect 168932 64268 168984 64320
rect 270500 64268 270552 64320
rect 69388 64200 69440 64252
rect 167644 64200 167696 64252
rect 169300 64200 169352 64252
rect 285680 64200 285732 64252
rect 168104 64132 168156 64184
rect 320180 64132 320232 64184
rect 110328 64064 110380 64116
rect 196624 64064 196676 64116
rect 166080 63588 166132 63640
rect 170404 63588 170456 63640
rect 167460 63520 167512 63572
rect 169944 63520 169996 63572
rect 169576 62908 169628 62960
rect 262220 62908 262272 62960
rect 167000 62840 167052 62892
rect 288440 62840 288492 62892
rect 169024 62772 169076 62824
rect 327080 62772 327132 62824
rect 169852 61480 169904 61532
rect 242900 61480 242952 61532
rect 169392 61412 169444 61464
rect 259552 61412 259604 61464
rect 167828 61344 167880 61396
rect 307024 61344 307076 61396
rect 203616 60664 203668 60716
rect 580172 60664 580224 60716
rect 168196 60052 168248 60104
rect 248420 60052 248472 60104
rect 169944 59984 169996 60036
rect 291200 59984 291252 60036
rect 196624 58624 196676 58676
rect 284300 58624 284352 58676
rect 169208 57196 169260 57248
rect 273260 57196 273312 57248
rect 170496 55904 170548 55956
rect 264244 55904 264296 55956
rect 169116 55836 169168 55888
rect 298100 55836 298152 55888
rect 194416 51688 194468 51740
rect 333980 51688 334032 51740
rect 168288 50328 168340 50380
rect 251272 50328 251324 50380
rect 178040 49036 178092 49088
rect 245660 49036 245712 49088
rect 169484 48968 169536 49020
rect 281540 48968 281592 49020
rect 171876 47540 171928 47592
rect 345020 47540 345072 47592
rect 164884 46860 164936 46912
rect 580172 46860 580224 46912
rect 186964 46180 187016 46232
rect 247040 46180 247092 46232
rect 2780 45500 2832 45552
rect 4804 45500 4856 45552
rect 170404 44820 170456 44872
rect 292672 44820 292724 44872
rect 167736 42032 167788 42084
rect 310520 42032 310572 42084
rect 167644 39312 167696 39364
rect 269120 39312 269172 39364
rect 194508 37884 194560 37936
rect 287060 37884 287112 37936
rect 171784 33736 171836 33788
rect 311164 33736 311216 33788
rect 2872 33056 2924 33108
rect 65524 33056 65576 33108
rect 191104 33056 191156 33108
rect 580172 33056 580224 33108
rect 190368 31016 190420 31068
rect 322940 31016 322992 31068
rect 167276 28228 167328 28280
rect 280160 28228 280212 28280
rect 169760 24080 169812 24132
rect 263600 24080 263652 24132
rect 220084 22720 220136 22772
rect 316132 22720 316184 22772
rect 198648 21360 198700 21412
rect 266360 21360 266412 21412
rect 3516 20612 3568 20664
rect 106372 20612 106424 20664
rect 188344 18572 188396 18624
rect 278780 18572 278832 18624
rect 209044 17212 209096 17264
rect 276020 17212 276072 17264
rect 169668 15852 169720 15904
rect 301504 15852 301556 15904
rect 173164 14424 173216 14476
rect 258264 14424 258316 14476
rect 167920 13064 167972 13116
rect 284392 13064 284444 13116
rect 175924 11704 175976 11756
rect 240140 11704 240192 11756
rect 259460 11704 259512 11756
rect 260656 11704 260708 11756
rect 185584 7624 185636 7676
rect 242992 7624 243044 7676
rect 206284 7556 206336 7608
rect 277124 7556 277176 7608
rect 182824 6808 182876 6860
rect 580172 6808 580224 6860
rect 187608 4972 187660 5024
rect 274824 4972 274876 5024
rect 180064 4904 180116 4956
rect 322112 4904 322164 4956
rect 181444 4836 181496 4888
rect 324412 4836 324464 4888
rect 4160 4768 4212 4820
rect 107660 4768 107712 4820
rect 174544 4768 174596 4820
rect 343364 4768 343416 4820
rect 235264 3680 235316 3732
rect 177396 3612 177448 3664
rect 245200 3748 245252 3800
rect 267740 3680 267792 3732
rect 242900 3612 242952 3664
rect 244096 3612 244148 3664
rect 251180 3612 251232 3664
rect 252376 3612 252428 3664
rect 284300 3612 284352 3664
rect 285036 3612 285088 3664
rect 299572 3612 299624 3664
rect 300768 3612 300820 3664
rect 311164 3612 311216 3664
rect 312636 3612 312688 3664
rect 203524 3544 203576 3596
rect 319720 3544 319772 3596
rect 324320 3544 324372 3596
rect 325608 3544 325660 3596
rect 332692 3544 332744 3596
rect 333888 3544 333940 3596
rect 184204 3476 184256 3528
rect 344560 3544 344612 3596
rect 340972 3476 341024 3528
rect 342168 3476 342220 3528
rect 349160 3476 349212 3528
rect 350448 3476 350500 3528
rect 69112 3408 69164 3460
rect 136456 3408 136508 3460
rect 177304 3408 177356 3460
rect 307024 3340 307076 3392
rect 309048 3340 309100 3392
rect 316040 3340 316092 3392
rect 317328 3340 317380 3392
rect 340972 3340 341024 3392
rect 264244 3136 264296 3188
rect 265348 3136 265400 3188
rect 572 2796 624 2848
rect 4160 2796 4212 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 8128 700330 8156 703520
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 24320 699718 24348 703520
rect 40512 700466 40540 703520
rect 40500 700460 40552 700466
rect 40500 700402 40552 700408
rect 72988 699718 73016 703520
rect 89180 700466 89208 703520
rect 78680 700460 78732 700466
rect 78680 700402 78732 700408
rect 89168 700460 89220 700466
rect 89168 700402 89220 700408
rect 73068 700392 73120 700398
rect 73068 700334 73120 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 25504 699712 25556 699718
rect 25504 699654 25556 699660
rect 66168 699712 66220 699718
rect 66168 699654 66220 699660
rect 72976 699712 73028 699718
rect 72976 699654 73028 699660
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 11704 565888 11756 565894
rect 11704 565830 11756 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 3424 514762 3476 514768
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 2778 475688 2834 475697
rect 2778 475623 2834 475632
rect 2792 474842 2820 475623
rect 2780 474836 2832 474842
rect 2780 474778 2832 474784
rect 4804 474836 4856 474842
rect 4804 474778 4856 474784
rect 3238 462632 3294 462641
rect 3238 462567 3294 462576
rect 3252 462398 3280 462567
rect 3240 462392 3292 462398
rect 3240 462334 3292 462340
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3436 422346 3464 423535
rect 3424 422340 3476 422346
rect 3424 422282 3476 422288
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3344 318850 3372 319223
rect 3332 318844 3384 318850
rect 3332 318786 3384 318792
rect 3330 293176 3386 293185
rect 3330 293111 3386 293120
rect 3344 292602 3372 293111
rect 3332 292596 3384 292602
rect 3332 292538 3384 292544
rect 3436 267734 3464 410479
rect 3516 397520 3568 397526
rect 3514 397488 3516 397497
rect 3568 397488 3570 397497
rect 3514 397423 3570 397432
rect 3606 371376 3662 371385
rect 3606 371311 3662 371320
rect 3514 358456 3570 358465
rect 3514 358391 3570 358400
rect 3344 267706 3464 267734
rect 3344 258738 3372 267706
rect 3422 267200 3478 267209
rect 3422 267135 3478 267144
rect 3436 266422 3464 267135
rect 3424 266416 3476 266422
rect 3424 266358 3476 266364
rect 3332 258732 3384 258738
rect 3332 258674 3384 258680
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3160 253978 3188 254079
rect 3148 253972 3200 253978
rect 3148 253914 3200 253920
rect 3054 241088 3110 241097
rect 3054 241023 3110 241032
rect 3068 240174 3096 241023
rect 3056 240168 3108 240174
rect 3056 240110 3108 240116
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3528 206281 3556 358391
rect 3620 260166 3648 371311
rect 3698 306232 3754 306241
rect 3698 306167 3754 306176
rect 3608 260160 3660 260166
rect 3608 260102 3660 260108
rect 3712 229094 3740 306167
rect 3712 229066 3832 229094
rect 3804 214606 3832 229066
rect 3792 214600 3844 214606
rect 3792 214542 3844 214548
rect 3514 206272 3570 206281
rect 3514 206207 3570 206216
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 3436 201550 3464 201855
rect 3424 201544 3476 201550
rect 3424 201486 3476 201492
rect 4816 200122 4844 474778
rect 10324 397520 10376 397526
rect 10324 397462 10376 397468
rect 7564 266416 7616 266422
rect 7564 266358 7616 266364
rect 4804 200116 4856 200122
rect 4804 200058 4856 200064
rect 7576 200054 7604 266358
rect 10336 256018 10364 397462
rect 10324 256012 10376 256018
rect 10324 255954 10376 255960
rect 10324 253972 10376 253978
rect 10324 253914 10376 253920
rect 10336 247722 10364 253914
rect 10324 247716 10376 247722
rect 10324 247658 10376 247664
rect 11716 205630 11744 565830
rect 18604 462392 18656 462398
rect 18604 462334 18656 462340
rect 15844 318844 15896 318850
rect 15844 318786 15896 318792
rect 15856 244934 15884 318786
rect 15844 244928 15896 244934
rect 15844 244870 15896 244876
rect 15844 225004 15896 225010
rect 15844 224946 15896 224952
rect 15856 215286 15884 224946
rect 15844 215280 15896 215286
rect 15844 215222 15896 215228
rect 11704 205624 11756 205630
rect 11704 205566 11756 205572
rect 7564 200048 7616 200054
rect 7564 199990 7616 199996
rect 18616 198626 18644 462334
rect 25516 257378 25544 699654
rect 55864 670744 55916 670750
rect 55864 670686 55916 670692
rect 54484 632120 54536 632126
rect 54484 632062 54536 632068
rect 25504 257372 25556 257378
rect 25504 257314 25556 257320
rect 54496 198665 54524 632062
rect 54482 198656 54538 198665
rect 18604 198620 18656 198626
rect 54482 198591 54538 198600
rect 18604 198562 18656 198568
rect 55876 198490 55904 670686
rect 62764 605872 62816 605878
rect 62764 605814 62816 605820
rect 61384 448588 61436 448594
rect 61384 448530 61436 448536
rect 58624 292596 58676 292602
rect 58624 292538 58676 292544
rect 58636 198558 58664 292538
rect 61396 199782 61424 448530
rect 62028 251592 62080 251598
rect 62028 251534 62080 251540
rect 61752 251388 61804 251394
rect 61752 251330 61804 251336
rect 61384 199776 61436 199782
rect 61384 199718 61436 199724
rect 58624 198552 58676 198558
rect 58624 198494 58676 198500
rect 55864 198484 55916 198490
rect 55864 198426 55916 198432
rect 3424 194608 3476 194614
rect 3424 194550 3476 194556
rect 3436 188873 3464 194550
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3422 162888 3478 162897
rect 3422 162823 3478 162832
rect 2962 149832 3018 149841
rect 2962 149767 3018 149776
rect 2976 149122 3004 149767
rect 2964 149116 3016 149122
rect 2964 149058 3016 149064
rect 3436 123486 3464 162823
rect 61764 137970 61792 251330
rect 61936 251252 61988 251258
rect 61936 251194 61988 251200
rect 61844 198076 61896 198082
rect 61844 198018 61896 198024
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 61752 137964 61804 137970
rect 61752 137906 61804 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3424 123480 3476 123486
rect 3424 123422 3476 123428
rect 60740 114504 60792 114510
rect 60740 114446 60792 114452
rect 60752 113830 60780 114446
rect 3516 113824 3568 113830
rect 3516 113766 3568 113772
rect 60740 113824 60792 113830
rect 60740 113766 60792 113772
rect 3424 111852 3476 111858
rect 3424 111794 3476 111800
rect 3436 110673 3464 111794
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3424 87032 3476 87038
rect 3424 86974 3476 86980
rect 3332 84856 3384 84862
rect 3332 84798 3384 84804
rect 3344 84194 3372 84798
rect 3436 84697 3464 86974
rect 3422 84688 3478 84697
rect 3422 84623 3478 84632
rect 3344 84166 3464 84194
rect 2870 71632 2926 71641
rect 2870 71567 2926 71576
rect 2884 67318 2912 71567
rect 2872 67312 2924 67318
rect 2872 67254 2924 67260
rect 2780 45552 2832 45558
rect 2778 45520 2780 45529
rect 2832 45520 2834 45529
rect 2778 45455 2834 45464
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2884 32473 2912 33050
rect 2870 32464 2926 32473
rect 2870 32399 2926 32408
rect 3436 6497 3464 84166
rect 3528 58585 3556 113766
rect 3606 97608 3662 97617
rect 3606 97543 3662 97552
rect 3620 70378 3648 97543
rect 4804 78736 4856 78742
rect 4804 78678 4856 78684
rect 3608 70372 3660 70378
rect 3608 70314 3660 70320
rect 3514 58576 3570 58585
rect 3514 58511 3570 58520
rect 4816 45558 4844 78678
rect 61856 68882 61884 198018
rect 61948 114374 61976 251194
rect 62040 114510 62068 251534
rect 62776 199850 62804 605814
rect 65524 579692 65576 579698
rect 65524 579634 65576 579640
rect 63408 251524 63460 251530
rect 63408 251466 63460 251472
rect 63316 250028 63368 250034
rect 63316 249970 63368 249976
rect 62764 199844 62816 199850
rect 62764 199786 62816 199792
rect 63224 198144 63276 198150
rect 63224 198086 63276 198092
rect 62028 114504 62080 114510
rect 62028 114446 62080 114452
rect 61936 114368 61988 114374
rect 61936 114310 61988 114316
rect 63236 68950 63264 198086
rect 63328 117298 63356 249970
rect 63316 117292 63368 117298
rect 63316 117234 63368 117240
rect 63420 111790 63448 251466
rect 64694 251424 64750 251433
rect 64694 251359 64750 251368
rect 64512 244928 64564 244934
rect 64512 244870 64564 244876
rect 64524 244322 64552 244870
rect 64512 244316 64564 244322
rect 64512 244258 64564 244264
rect 63500 225616 63552 225622
rect 63500 225558 63552 225564
rect 63512 225010 63540 225558
rect 63500 225004 63552 225010
rect 63500 224946 63552 224952
rect 64420 215348 64472 215354
rect 64420 215290 64472 215296
rect 63500 201544 63552 201550
rect 63500 201486 63552 201492
rect 63512 193866 63540 201486
rect 63500 193860 63552 193866
rect 63500 193802 63552 193808
rect 64432 189786 64460 215290
rect 64524 199918 64552 244258
rect 64604 225616 64656 225622
rect 64604 225558 64656 225564
rect 64512 199912 64564 199918
rect 64512 199854 64564 199860
rect 64420 189780 64472 189786
rect 64420 189722 64472 189728
rect 64420 116068 64472 116074
rect 64420 116010 64472 116016
rect 64328 115116 64380 115122
rect 64328 115058 64380 115064
rect 64236 114776 64288 114782
rect 64236 114718 64288 114724
rect 63408 111784 63460 111790
rect 63408 111726 63460 111732
rect 64248 96626 64276 114718
rect 64340 99346 64368 115058
rect 64328 99340 64380 99346
rect 64328 99282 64380 99288
rect 64236 96620 64288 96626
rect 64236 96562 64288 96568
rect 64432 92478 64460 116010
rect 64524 113286 64552 199854
rect 64616 113830 64644 225558
rect 64708 118658 64736 251359
rect 64788 249824 64840 249830
rect 64788 249766 64840 249772
rect 64696 118652 64748 118658
rect 64696 118594 64748 118600
rect 64800 117230 64828 249766
rect 65338 210216 65394 210225
rect 65338 210151 65394 210160
rect 64788 117224 64840 117230
rect 64788 117166 64840 117172
rect 64696 116000 64748 116006
rect 64696 115942 64748 115948
rect 64604 113824 64656 113830
rect 64604 113766 64656 113772
rect 64512 113280 64564 113286
rect 64512 113222 64564 113228
rect 64524 104854 64552 113222
rect 64512 104848 64564 104854
rect 64512 104790 64564 104796
rect 64708 93838 64736 115942
rect 64788 114572 64840 114578
rect 64788 114514 64840 114520
rect 64800 103494 64828 114514
rect 64788 103488 64840 103494
rect 64788 103430 64840 103436
rect 64696 93832 64748 93838
rect 64696 93774 64748 93780
rect 64420 92472 64472 92478
rect 64420 92414 64472 92420
rect 65352 78606 65380 210151
rect 65430 200288 65486 200297
rect 65430 200223 65486 200232
rect 65444 78674 65472 200223
rect 65536 199714 65564 579634
rect 65892 254788 65944 254794
rect 65892 254730 65944 254736
rect 65800 230512 65852 230518
rect 65800 230454 65852 230460
rect 65616 220856 65668 220862
rect 65616 220798 65668 220804
rect 65524 199708 65576 199714
rect 65524 199650 65576 199656
rect 65628 199442 65656 220798
rect 65708 204332 65760 204338
rect 65708 204274 65760 204280
rect 65616 199436 65668 199442
rect 65616 199378 65668 199384
rect 65720 175982 65748 204274
rect 65812 199170 65840 230454
rect 65904 230450 65932 254730
rect 66076 251660 66128 251666
rect 66076 251602 66128 251608
rect 65982 251560 66038 251569
rect 65982 251495 66038 251504
rect 65892 230444 65944 230450
rect 65892 230386 65944 230392
rect 65892 218068 65944 218074
rect 65892 218010 65944 218016
rect 65800 199164 65852 199170
rect 65800 199106 65852 199112
rect 65800 198212 65852 198218
rect 65800 198154 65852 198160
rect 65708 175976 65760 175982
rect 65708 175918 65760 175924
rect 65524 137964 65576 137970
rect 65524 137906 65576 137912
rect 65536 114442 65564 137906
rect 65708 114640 65760 114646
rect 65708 114582 65760 114588
rect 65524 114436 65576 114442
rect 65524 114378 65576 114384
rect 65524 112056 65576 112062
rect 65524 111998 65576 112004
rect 65432 78668 65484 78674
rect 65432 78610 65484 78616
rect 65340 78600 65392 78606
rect 65340 78542 65392 78548
rect 63224 68944 63276 68950
rect 63224 68886 63276 68892
rect 61844 68876 61896 68882
rect 61844 68818 61896 68824
rect 4804 45552 4856 45558
rect 4804 45494 4856 45500
rect 65536 33114 65564 111998
rect 65720 92410 65748 114582
rect 65708 92404 65760 92410
rect 65708 92346 65760 92352
rect 65812 68746 65840 198154
rect 65904 198014 65932 218010
rect 65892 198008 65944 198014
rect 65892 197950 65944 197956
rect 65996 118590 66024 251495
rect 65984 118584 66036 118590
rect 65984 118526 66036 118532
rect 65984 117360 66036 117366
rect 65984 117302 66036 117308
rect 65996 97986 66024 117302
rect 66088 114238 66116 251602
rect 66180 198422 66208 699654
rect 71780 345092 71832 345098
rect 71780 345034 71832 345040
rect 68744 254584 68796 254590
rect 68744 254526 68796 254532
rect 67548 254448 67600 254454
rect 67548 254390 67600 254396
rect 67456 254176 67508 254182
rect 67456 254118 67508 254124
rect 67088 249144 67140 249150
rect 67088 249086 67140 249092
rect 66996 243500 67048 243506
rect 66996 243442 67048 243448
rect 66904 240168 66956 240174
rect 66904 240110 66956 240116
rect 66628 232620 66680 232626
rect 66628 232562 66680 232568
rect 66168 198416 66220 198422
rect 66168 198358 66220 198364
rect 66168 114844 66220 114850
rect 66168 114786 66220 114792
rect 66076 114232 66128 114238
rect 66076 114174 66128 114180
rect 66074 112160 66130 112169
rect 66074 112095 66130 112104
rect 66088 100706 66116 112095
rect 66076 100700 66128 100706
rect 66076 100642 66128 100648
rect 66180 100638 66208 114786
rect 66168 100632 66220 100638
rect 66168 100574 66220 100580
rect 65984 97980 66036 97986
rect 65984 97922 66036 97928
rect 66640 96558 66668 232562
rect 66916 225350 66944 240110
rect 66904 225344 66956 225350
rect 66904 225286 66956 225292
rect 66902 223816 66958 223825
rect 66902 223751 66958 223760
rect 66812 216708 66864 216714
rect 66812 216650 66864 216656
rect 66720 201544 66772 201550
rect 66720 201486 66772 201492
rect 66732 173194 66760 201486
rect 66824 191146 66852 216650
rect 66916 197985 66944 223751
rect 66902 197976 66958 197985
rect 66902 197911 66958 197920
rect 66812 191140 66864 191146
rect 66812 191082 66864 191088
rect 66720 173188 66772 173194
rect 66720 173130 66772 173136
rect 66628 96552 66680 96558
rect 66628 96494 66680 96500
rect 65984 78736 66036 78742
rect 65984 78678 66036 78684
rect 65996 69902 66024 78678
rect 66168 78668 66220 78674
rect 66168 78610 66220 78616
rect 66076 78600 66128 78606
rect 66076 78542 66128 78548
rect 65984 69896 66036 69902
rect 65984 69838 66036 69844
rect 65800 68740 65852 68746
rect 65800 68682 65852 68688
rect 66088 64802 66116 78542
rect 66180 77654 66208 78610
rect 66168 77648 66220 77654
rect 66168 77590 66220 77596
rect 66180 64870 66208 77590
rect 66732 72486 66760 173130
rect 66824 83609 66852 191082
rect 66916 88534 66944 197911
rect 67008 126274 67036 243442
rect 67100 240990 67128 249086
rect 67468 241641 67496 254118
rect 67560 249150 67588 254390
rect 68756 253934 68784 254526
rect 69296 254380 69348 254386
rect 69296 254322 69348 254328
rect 69020 254312 69072 254318
rect 69020 254254 69072 254260
rect 68756 253906 68968 253934
rect 68468 253496 68520 253502
rect 68468 253438 68520 253444
rect 68284 253020 68336 253026
rect 68284 252962 68336 252968
rect 68192 250708 68244 250714
rect 68192 250650 68244 250656
rect 68008 250368 68060 250374
rect 68008 250310 68060 250316
rect 67916 250096 67968 250102
rect 67916 250038 67968 250044
rect 67548 249144 67600 249150
rect 67548 249086 67600 249092
rect 67638 247752 67694 247761
rect 67638 247687 67640 247696
rect 67692 247687 67694 247696
rect 67640 247658 67692 247664
rect 67546 245576 67602 245585
rect 67546 245511 67602 245520
rect 67454 241632 67510 241641
rect 67454 241567 67510 241576
rect 67088 240984 67140 240990
rect 67088 240926 67140 240932
rect 66996 126268 67048 126274
rect 66996 126210 67048 126216
rect 67008 104145 67036 126210
rect 67100 112130 67128 240926
rect 67560 238754 67588 245511
rect 67638 244352 67694 244361
rect 67638 244287 67640 244296
rect 67692 244287 67694 244296
rect 67640 244258 67692 244264
rect 67284 238726 67588 238754
rect 67928 238754 67956 250038
rect 68020 243250 68048 250310
rect 68204 243642 68232 250650
rect 68296 245585 68324 252962
rect 68376 249960 68428 249966
rect 68376 249902 68428 249908
rect 68282 245576 68338 245585
rect 68282 245511 68338 245520
rect 68192 243636 68244 243642
rect 68192 243578 68244 243584
rect 68388 243574 68416 249902
rect 68376 243568 68428 243574
rect 68376 243510 68428 243516
rect 68020 243222 68324 243250
rect 68296 238754 68324 243222
rect 68376 240984 68428 240990
rect 68374 240952 68376 240961
rect 68428 240952 68430 240961
rect 68374 240887 68430 240896
rect 67928 238726 68232 238754
rect 68296 238726 68416 238754
rect 67180 200184 67232 200190
rect 67180 200126 67232 200132
rect 67088 112124 67140 112130
rect 67088 112066 67140 112072
rect 67100 111926 67128 112066
rect 67088 111920 67140 111926
rect 67088 111862 67140 111868
rect 66994 104136 67050 104145
rect 66994 104071 67050 104080
rect 66904 88528 66956 88534
rect 66904 88470 66956 88476
rect 66810 83600 66866 83609
rect 66810 83535 66866 83544
rect 67192 74534 67220 200126
rect 67284 114306 67312 238726
rect 67638 230616 67694 230625
rect 67638 230551 67694 230560
rect 67652 230518 67680 230551
rect 67640 230512 67692 230518
rect 67640 230454 67692 230460
rect 67732 230444 67784 230450
rect 67732 230386 67784 230392
rect 67744 229401 67772 230386
rect 67730 229392 67786 229401
rect 67730 229327 67786 229336
rect 68204 225865 68232 238726
rect 68388 236881 68416 238726
rect 68374 236872 68430 236881
rect 68374 236807 68430 236816
rect 68480 235362 68508 253438
rect 68744 253156 68796 253162
rect 68744 253098 68796 253104
rect 68652 250300 68704 250306
rect 68652 250242 68704 250248
rect 68558 247752 68614 247761
rect 68558 247687 68614 247696
rect 68388 235334 68508 235362
rect 68388 232121 68416 235334
rect 68468 233912 68520 233918
rect 68468 233854 68520 233860
rect 68374 232112 68430 232121
rect 68374 232047 68430 232056
rect 68480 228041 68508 233854
rect 68466 228032 68522 228041
rect 68466 227967 68522 227976
rect 67822 225856 67878 225865
rect 67822 225791 67878 225800
rect 68190 225856 68246 225865
rect 68190 225791 68246 225800
rect 67836 225622 67864 225791
rect 67824 225616 67876 225622
rect 67824 225558 67876 225564
rect 68006 221096 68062 221105
rect 68006 221031 68062 221040
rect 68020 220862 68048 221031
rect 68008 220856 68060 220862
rect 68008 220798 68060 220804
rect 67456 219496 67508 219502
rect 67456 219438 67508 219444
rect 67364 205692 67416 205698
rect 67364 205634 67416 205640
rect 67272 114300 67324 114306
rect 67272 114242 67324 114248
rect 67272 111920 67324 111926
rect 67272 111862 67324 111868
rect 67284 101425 67312 111862
rect 67270 101416 67326 101425
rect 67270 101351 67326 101360
rect 67376 82414 67404 205634
rect 67468 86970 67496 219438
rect 68190 219056 68246 219065
rect 68190 218991 68246 219000
rect 68204 218074 68232 218991
rect 68466 218376 68522 218385
rect 68466 218311 68522 218320
rect 68192 218068 68244 218074
rect 68192 218010 68244 218016
rect 68374 217016 68430 217025
rect 68374 216951 68430 216960
rect 68388 216714 68416 216951
rect 68376 216708 68428 216714
rect 68376 216650 68428 216656
rect 67638 216336 67694 216345
rect 67638 216271 67694 216280
rect 67652 215354 67680 216271
rect 67640 215348 67692 215354
rect 67640 215290 67692 215296
rect 68374 214976 68430 214985
rect 68374 214911 68430 214920
rect 67640 214600 67692 214606
rect 67640 214542 67692 214548
rect 67652 214441 67680 214542
rect 67638 214432 67694 214441
rect 67638 214367 67694 214376
rect 68190 214432 68246 214441
rect 68190 214367 68246 214376
rect 67914 213616 67970 213625
rect 67914 213551 67970 213560
rect 67730 206272 67786 206281
rect 67730 206207 67786 206216
rect 67638 202736 67694 202745
rect 67638 202671 67694 202680
rect 67652 201550 67680 202671
rect 67640 201544 67692 201550
rect 67640 201486 67692 201492
rect 67744 180985 67772 206207
rect 67824 205624 67876 205630
rect 67822 205592 67824 205601
rect 67876 205592 67878 205601
rect 67822 205527 67878 205536
rect 67928 199374 67956 213551
rect 68008 204944 68060 204950
rect 68008 204886 68060 204892
rect 67916 199368 67968 199374
rect 67916 199310 67968 199316
rect 68020 184890 68048 204886
rect 68098 204776 68154 204785
rect 68098 204711 68154 204720
rect 68112 204338 68140 204711
rect 68100 204332 68152 204338
rect 68100 204274 68152 204280
rect 68204 186697 68232 214367
rect 68388 205698 68416 214911
rect 68376 205692 68428 205698
rect 68376 205634 68428 205640
rect 68388 201249 68416 205634
rect 68374 201240 68430 201249
rect 68374 201175 68430 201184
rect 68480 192506 68508 218311
rect 68572 198694 68600 247687
rect 68664 243681 68692 250242
rect 68756 249801 68784 253098
rect 68836 250232 68888 250238
rect 68836 250174 68888 250180
rect 68742 249792 68798 249801
rect 68742 249727 68798 249736
rect 68744 248600 68796 248606
rect 68744 248542 68796 248548
rect 68650 243672 68706 243681
rect 68650 243607 68706 243616
rect 68652 243568 68704 243574
rect 68652 243510 68704 243516
rect 68664 230081 68692 243510
rect 68756 233918 68784 248542
rect 68848 248305 68876 250174
rect 68834 248296 68890 248305
rect 68834 248231 68890 248240
rect 68836 243636 68888 243642
rect 68836 243578 68888 243584
rect 68848 237561 68876 243578
rect 68834 237552 68890 237561
rect 68834 237487 68890 237496
rect 68744 233912 68796 233918
rect 68744 233854 68796 233860
rect 68742 232656 68798 232665
rect 68742 232591 68744 232600
rect 68796 232591 68798 232600
rect 68744 232562 68796 232568
rect 68650 230072 68706 230081
rect 68650 230007 68706 230016
rect 68940 227361 68968 253906
rect 69032 234161 69060 254254
rect 69204 252068 69256 252074
rect 69204 252010 69256 252016
rect 69110 246256 69166 246265
rect 69110 246191 69166 246200
rect 69018 234152 69074 234161
rect 69018 234087 69074 234096
rect 68926 227352 68982 227361
rect 68926 227287 68982 227296
rect 68744 225344 68796 225350
rect 68742 225312 68744 225321
rect 68796 225312 68798 225321
rect 68742 225247 68798 225256
rect 69018 225312 69074 225321
rect 69018 225247 69074 225256
rect 68650 223136 68706 223145
rect 68650 223071 68706 223080
rect 68664 215294 68692 223071
rect 68926 220416 68982 220425
rect 68926 220351 68982 220360
rect 68940 219502 68968 220351
rect 68928 219496 68980 219502
rect 68928 219438 68980 219444
rect 68664 215266 68784 215294
rect 68650 201376 68706 201385
rect 68650 201311 68706 201320
rect 68560 198688 68612 198694
rect 68560 198630 68612 198636
rect 68468 192500 68520 192506
rect 68468 192442 68520 192448
rect 68190 186688 68246 186697
rect 68190 186623 68246 186632
rect 68008 184884 68060 184890
rect 68008 184826 68060 184832
rect 67730 180976 67786 180985
rect 67730 180911 67786 180920
rect 67548 114300 67600 114306
rect 67548 114242 67600 114248
rect 67560 113558 67588 114242
rect 67548 113552 67600 113558
rect 67548 113494 67600 113500
rect 67560 105505 67588 113494
rect 67546 105496 67602 105505
rect 67546 105431 67602 105440
rect 67640 104848 67692 104854
rect 67638 104816 67640 104825
rect 67692 104816 67694 104825
rect 67638 104751 67694 104760
rect 67640 103488 67692 103494
rect 67640 103430 67692 103436
rect 67652 102785 67680 103430
rect 67638 102776 67694 102785
rect 67638 102711 67694 102720
rect 67638 100736 67694 100745
rect 67638 100671 67640 100680
rect 67692 100671 67694 100680
rect 67640 100642 67692 100648
rect 67640 99340 67692 99346
rect 67640 99282 67692 99288
rect 67652 98705 67680 99282
rect 67638 98696 67694 98705
rect 67638 98631 67694 98640
rect 67640 97980 67692 97986
rect 67640 97922 67692 97928
rect 67652 97889 67680 97922
rect 67638 97880 67694 97889
rect 67638 97815 67694 97824
rect 67640 96620 67692 96626
rect 67640 96562 67692 96568
rect 67652 95985 67680 96562
rect 67638 95976 67694 95985
rect 67638 95911 67694 95920
rect 67640 93832 67692 93838
rect 67640 93774 67692 93780
rect 67652 93265 67680 93774
rect 67638 93256 67694 93265
rect 67638 93191 67694 93200
rect 67640 92472 67692 92478
rect 67640 92414 67692 92420
rect 67652 91225 67680 92414
rect 67638 91216 67694 91225
rect 67638 91151 67694 91160
rect 67456 86964 67508 86970
rect 67456 86906 67508 86912
rect 67640 84856 67692 84862
rect 67640 84798 67692 84804
rect 67652 84425 67680 84798
rect 67638 84416 67694 84425
rect 67638 84351 67694 84360
rect 67364 82408 67416 82414
rect 67364 82350 67416 82356
rect 67638 78840 67694 78849
rect 67638 78775 67694 78784
rect 67652 78742 67680 78775
rect 67640 78736 67692 78742
rect 67640 78678 67692 78684
rect 67640 78600 67692 78606
rect 67640 78542 67692 78548
rect 67652 78305 67680 78542
rect 67638 78296 67694 78305
rect 67638 78231 67694 78240
rect 67640 77648 67692 77654
rect 67638 77616 67640 77625
rect 67692 77616 67694 77625
rect 67638 77551 67694 77560
rect 67744 75857 67772 180911
rect 67916 112396 67968 112402
rect 67916 112338 67968 112344
rect 67824 111920 67876 111926
rect 67824 111862 67876 111868
rect 67836 84862 67864 111862
rect 67928 87825 67956 112338
rect 67914 87816 67970 87825
rect 67914 87751 67970 87760
rect 67916 86964 67968 86970
rect 67916 86906 67968 86912
rect 67928 85785 67956 86906
rect 67914 85776 67970 85785
rect 67914 85711 67970 85720
rect 67824 84856 67876 84862
rect 67824 84798 67876 84804
rect 67822 80880 67878 80889
rect 67822 80815 67878 80824
rect 67730 75848 67786 75857
rect 67730 75783 67786 75792
rect 67192 74506 67588 74534
rect 66720 72480 66772 72486
rect 66720 72422 66772 72428
rect 67560 70106 67588 74506
rect 67548 70100 67600 70106
rect 67548 70042 67600 70048
rect 66168 64864 66220 64870
rect 66168 64806 66220 64812
rect 66076 64796 66128 64802
rect 66076 64738 66128 64744
rect 67560 64734 67588 70042
rect 67836 66774 67864 80815
rect 67824 66768 67876 66774
rect 67824 66710 67876 66716
rect 67928 65958 67956 85711
rect 68020 78849 68048 184826
rect 68100 92404 68152 92410
rect 68100 92346 68152 92352
rect 68112 91905 68140 92346
rect 68098 91896 68154 91905
rect 68098 91831 68154 91840
rect 68100 87032 68152 87038
rect 68098 87000 68100 87009
rect 68152 87000 68154 87009
rect 68098 86935 68154 86944
rect 68204 80889 68232 186623
rect 68480 112198 68508 192442
rect 68572 113354 68600 198630
rect 68664 172514 68692 201311
rect 68756 199578 68784 215266
rect 68834 208176 68890 208185
rect 68834 208111 68890 208120
rect 68744 199572 68796 199578
rect 68744 199514 68796 199520
rect 68848 198762 68876 208111
rect 68940 204921 68968 219438
rect 68926 204912 68982 204921
rect 68926 204847 68982 204856
rect 69032 199510 69060 225247
rect 69020 199504 69072 199510
rect 69020 199446 69072 199452
rect 68836 198756 68888 198762
rect 68836 198698 68888 198704
rect 68928 177336 68980 177342
rect 68926 177304 68928 177313
rect 68980 177304 68982 177313
rect 68926 177239 68982 177248
rect 68652 172508 68704 172514
rect 68652 172450 68704 172456
rect 68560 113348 68612 113354
rect 68560 113290 68612 113296
rect 68468 112192 68520 112198
rect 68468 112134 68520 112140
rect 68480 111926 68508 112134
rect 68468 111920 68520 111926
rect 68468 111862 68520 111868
rect 68572 106865 68600 113290
rect 68558 106856 68614 106865
rect 68558 106791 68614 106800
rect 68284 100632 68336 100638
rect 68284 100574 68336 100580
rect 68296 100065 68324 100574
rect 68282 100056 68338 100065
rect 68282 99991 68338 100000
rect 68558 89040 68614 89049
rect 68558 88975 68614 88984
rect 68468 88528 68520 88534
rect 68466 88496 68468 88505
rect 68520 88496 68522 88505
rect 68466 88431 68522 88440
rect 68480 84194 68508 88431
rect 68388 84166 68508 84194
rect 68190 80880 68246 80889
rect 68190 80815 68246 80824
rect 68006 78840 68062 78849
rect 68006 78775 68062 78784
rect 68284 72480 68336 72486
rect 68284 72422 68336 72428
rect 68296 72049 68324 72422
rect 68282 72040 68338 72049
rect 68282 71975 68338 71984
rect 67916 65952 67968 65958
rect 67916 65894 67968 65900
rect 68296 65793 68324 71975
rect 68388 69698 68416 84166
rect 68468 82408 68520 82414
rect 68468 82350 68520 82356
rect 68480 81569 68508 82350
rect 68466 81560 68522 81569
rect 68466 81495 68522 81504
rect 68376 69692 68428 69698
rect 68376 69634 68428 69640
rect 68480 67289 68508 81495
rect 68572 69766 68600 88975
rect 68664 71369 68692 172450
rect 68834 117328 68890 117337
rect 68834 117263 68890 117272
rect 68848 116113 68876 117263
rect 68834 116104 68890 116113
rect 68834 116039 68890 116048
rect 68744 112328 68796 112334
rect 68744 112270 68796 112276
rect 68756 103514 68784 112270
rect 68848 107545 68876 116039
rect 68928 111920 68980 111926
rect 68928 111862 68980 111868
rect 68940 111790 68968 111862
rect 68928 111784 68980 111790
rect 68928 111726 68980 111732
rect 68834 107536 68890 107545
rect 68834 107471 68890 107480
rect 68756 103486 68968 103514
rect 68940 94625 68968 103486
rect 68926 94616 68982 94625
rect 68926 94551 68982 94560
rect 69032 89049 69060 199446
rect 69124 196722 69152 246191
rect 69112 196716 69164 196722
rect 69112 196658 69164 196664
rect 69216 111722 69244 252010
rect 69308 234841 69336 254322
rect 69388 254244 69440 254250
rect 69388 254186 69440 254192
rect 69400 236201 69428 254186
rect 69480 252748 69532 252754
rect 69480 252690 69532 252696
rect 69492 243545 69520 252690
rect 71792 252074 71820 345034
rect 71780 252068 71832 252074
rect 71780 252010 71832 252016
rect 72608 252068 72660 252074
rect 72608 252010 72660 252016
rect 71320 251932 71372 251938
rect 71320 251874 71372 251880
rect 71332 249764 71360 251874
rect 71962 251832 72018 251841
rect 71962 251767 72018 251776
rect 71976 249764 72004 251767
rect 72620 249764 72648 252010
rect 73080 251841 73108 700334
rect 75920 683188 75972 683194
rect 75920 683130 75972 683136
rect 73896 254108 73948 254114
rect 73896 254050 73948 254056
rect 73066 251832 73122 251841
rect 73066 251767 73122 251776
rect 73908 249764 73936 254050
rect 75828 251864 75880 251870
rect 75828 251806 75880 251812
rect 74540 251524 74592 251530
rect 74540 251466 74592 251472
rect 74552 249764 74580 251466
rect 75840 251258 75868 251806
rect 75932 251666 75960 683130
rect 77760 254040 77812 254046
rect 77760 253982 77812 253988
rect 75920 251660 75972 251666
rect 75920 251602 75972 251608
rect 76472 251660 76524 251666
rect 76472 251602 76524 251608
rect 75828 251252 75880 251258
rect 75828 251194 75880 251200
rect 75840 249764 75868 251194
rect 76484 249764 76512 251602
rect 77772 249764 77800 253982
rect 78402 249928 78458 249937
rect 78402 249863 78458 249872
rect 78416 249764 78444 249863
rect 78692 249830 78720 700402
rect 105464 700330 105492 703520
rect 122840 700460 122892 700466
rect 122840 700402 122892 700408
rect 94504 700324 94556 700330
rect 94504 700266 94556 700272
rect 105452 700324 105504 700330
rect 105452 700266 105504 700272
rect 120724 700324 120776 700330
rect 120724 700266 120776 700272
rect 94516 267734 94544 700266
rect 95884 656940 95936 656946
rect 95884 656882 95936 656888
rect 94516 267706 94728 267734
rect 91284 254652 91336 254658
rect 91284 254594 91336 254600
rect 80980 253564 81032 253570
rect 80980 253506 81032 253512
rect 80336 252136 80388 252142
rect 80336 252078 80388 252084
rect 78680 249824 78732 249830
rect 79232 249824 79284 249830
rect 78680 249766 78732 249772
rect 79074 249772 79232 249778
rect 79074 249766 79284 249772
rect 79074 249750 79272 249766
rect 80348 249764 80376 252078
rect 80992 251394 81020 253506
rect 85488 253224 85540 253230
rect 85488 253166 85540 253172
rect 85500 251598 85528 253166
rect 90640 252952 90692 252958
rect 90640 252894 90692 252900
rect 89352 252816 89404 252822
rect 89352 252758 89404 252764
rect 85488 251592 85540 251598
rect 84198 251560 84254 251569
rect 85488 251534 85540 251540
rect 86776 251592 86828 251598
rect 86776 251534 86828 251540
rect 84198 251495 84254 251504
rect 80980 251388 81032 251394
rect 80980 251330 81032 251336
rect 80992 249764 81020 251330
rect 82912 250436 82964 250442
rect 82912 250378 82964 250384
rect 82266 250064 82322 250073
rect 82924 250034 82952 250378
rect 82266 249999 82322 250008
rect 82912 250028 82964 250034
rect 82280 249764 82308 249999
rect 82912 249970 82964 249976
rect 82924 249764 82952 249970
rect 84212 249764 84240 251495
rect 84842 251424 84898 251433
rect 84842 251359 84898 251368
rect 84856 249764 84884 251359
rect 85500 249764 85528 251534
rect 86788 249764 86816 251534
rect 88706 250200 88762 250209
rect 88706 250135 88762 250144
rect 87420 250096 87472 250102
rect 87420 250038 87472 250044
rect 87432 249764 87460 250038
rect 88720 249764 88748 250135
rect 89364 249764 89392 252758
rect 90652 249764 90680 252894
rect 91296 249764 91324 254594
rect 91928 254516 91980 254522
rect 91928 254458 91980 254464
rect 91940 249764 91968 254458
rect 93216 253292 93268 253298
rect 93216 253234 93268 253240
rect 93228 249764 93256 253234
rect 93860 253088 93912 253094
rect 93860 253030 93912 253036
rect 93872 249764 93900 253030
rect 94700 251705 94728 267706
rect 94686 251696 94742 251705
rect 94686 251631 94742 251640
rect 95148 251660 95200 251666
rect 94700 249778 94728 251631
rect 95148 251602 95200 251608
rect 95160 250481 95188 251602
rect 95896 250578 95924 656882
rect 106280 618316 106332 618322
rect 106280 618258 106332 618264
rect 99380 501016 99432 501022
rect 99380 500958 99432 500964
rect 99012 253428 99064 253434
rect 99012 253370 99064 253376
rect 97080 251660 97132 251666
rect 97080 251602 97132 251608
rect 95884 250572 95936 250578
rect 95884 250514 95936 250520
rect 95146 250472 95202 250481
rect 95146 250407 95202 250416
rect 95896 249778 95924 250514
rect 94700 249750 95174 249778
rect 95818 249750 95924 249778
rect 97092 249764 97120 251602
rect 97724 251320 97776 251326
rect 97724 251262 97776 251268
rect 97736 249764 97764 251262
rect 99024 249764 99052 253370
rect 99392 249778 99420 500958
rect 104164 254720 104216 254726
rect 104164 254662 104216 254668
rect 103520 252612 103572 252618
rect 103520 252554 103572 252560
rect 102232 252000 102284 252006
rect 102232 251942 102284 251948
rect 101588 251728 101640 251734
rect 101588 251670 101640 251676
rect 100300 251252 100352 251258
rect 100300 251194 100352 251200
rect 99656 250028 99708 250034
rect 99656 249970 99708 249976
rect 99668 249778 99696 249970
rect 99392 249764 99696 249778
rect 100312 249764 100340 251194
rect 101600 249764 101628 251670
rect 102244 249764 102272 251942
rect 103428 251320 103480 251326
rect 103428 251262 103480 251268
rect 103440 251161 103468 251262
rect 103426 251152 103482 251161
rect 103426 251087 103482 251096
rect 103532 249764 103560 252554
rect 104176 249764 104204 254662
rect 105452 252204 105504 252210
rect 105452 252146 105504 252152
rect 105464 249764 105492 252146
rect 106094 251968 106150 251977
rect 106094 251903 106150 251912
rect 106108 249764 106136 251903
rect 106292 249778 106320 618258
rect 107660 514820 107712 514826
rect 107660 514762 107712 514768
rect 107672 251190 107700 514762
rect 119344 422340 119396 422346
rect 119344 422282 119396 422288
rect 119356 267734 119384 422282
rect 119356 267706 119476 267734
rect 114468 253972 114520 253978
rect 114468 253914 114520 253920
rect 111892 252884 111944 252890
rect 111892 252826 111944 252832
rect 109960 252272 110012 252278
rect 109960 252214 110012 252220
rect 108028 251796 108080 251802
rect 108028 251738 108080 251744
rect 107660 251184 107712 251190
rect 107660 251126 107712 251132
rect 106740 249892 106792 249898
rect 106740 249834 106792 249840
rect 106752 249778 106780 249834
rect 106292 249764 106780 249778
rect 108040 249764 108068 251738
rect 108672 251184 108724 251190
rect 108672 251126 108724 251132
rect 108684 250646 108712 251126
rect 108672 250640 108724 250646
rect 108672 250582 108724 250588
rect 108684 249764 108712 250582
rect 109972 249764 110000 252214
rect 110604 251388 110656 251394
rect 110604 251330 110656 251336
rect 110616 249764 110644 251330
rect 111904 249764 111932 252826
rect 112536 252680 112588 252686
rect 112536 252622 112588 252628
rect 112168 252136 112220 252142
rect 112168 252078 112220 252084
rect 112180 249801 112208 252078
rect 112166 249792 112222 249801
rect 99392 249750 99682 249764
rect 106292 249750 106766 249764
rect 112548 249764 112576 252622
rect 113180 252136 113232 252142
rect 113180 252078 113232 252084
rect 113192 249764 113220 252078
rect 114480 249764 114508 253914
rect 119158 252920 119214 252929
rect 119158 252855 119214 252864
rect 118056 252272 118108 252278
rect 118056 252214 118108 252220
rect 117044 251456 117096 251462
rect 117044 251398 117096 251404
rect 116398 251288 116454 251297
rect 116398 251223 116454 251232
rect 116412 249764 116440 251223
rect 117056 249764 117084 251398
rect 117228 251252 117280 251258
rect 117228 251194 117280 251200
rect 117240 250578 117268 251194
rect 117964 250776 118016 250782
rect 117964 250718 118016 250724
rect 117228 250572 117280 250578
rect 117228 250514 117280 250520
rect 117976 250238 118004 250718
rect 117964 250232 118016 250238
rect 117964 250174 118016 250180
rect 112166 249727 112222 249736
rect 115480 249552 115532 249558
rect 115138 249500 115480 249506
rect 115138 249494 115532 249500
rect 115138 249478 115520 249494
rect 118068 249490 118096 252214
rect 118792 252204 118844 252210
rect 118792 252146 118844 252152
rect 118698 251424 118754 251433
rect 118698 251359 118754 251368
rect 118332 251320 118384 251326
rect 118332 251262 118384 251268
rect 118344 249764 118372 251262
rect 118712 249762 118740 251359
rect 118700 249756 118752 249762
rect 118700 249698 118752 249704
rect 118804 249490 118832 252146
rect 118976 251252 119028 251258
rect 118976 251194 119028 251200
rect 118988 249764 119016 251194
rect 119172 249694 119200 252855
rect 119250 251696 119306 251705
rect 119250 251631 119306 251640
rect 119160 249688 119212 249694
rect 119160 249630 119212 249636
rect 119160 249552 119212 249558
rect 119160 249494 119212 249500
rect 118056 249484 118108 249490
rect 118056 249426 118108 249432
rect 118792 249484 118844 249490
rect 118792 249426 118844 249432
rect 69860 249206 70058 249234
rect 69860 248470 69888 249206
rect 119172 248538 119200 249494
rect 119160 248532 119212 248538
rect 119160 248474 119212 248480
rect 69848 248464 69900 248470
rect 69848 248406 69900 248412
rect 119264 247790 119292 251631
rect 119342 249928 119398 249937
rect 119342 249863 119398 249872
rect 119252 247784 119304 247790
rect 119252 247726 119304 247732
rect 69478 243536 69534 243545
rect 69478 243471 69480 243480
rect 69532 243471 69534 243480
rect 69480 243442 69532 243448
rect 69386 236192 69442 236201
rect 69386 236127 69442 236136
rect 69294 234832 69350 234841
rect 69294 234767 69350 234776
rect 119356 233102 119384 249863
rect 119448 249778 119476 267706
rect 120172 260160 120224 260166
rect 120172 260102 120224 260108
rect 119988 252612 120040 252618
rect 119988 252554 120040 252560
rect 119894 251832 119950 251841
rect 119894 251767 119950 251776
rect 119804 249824 119856 249830
rect 119448 249750 119752 249778
rect 119804 249766 119856 249772
rect 119436 249688 119488 249694
rect 119436 249630 119488 249636
rect 119344 233096 119396 233102
rect 119344 233038 119396 233044
rect 119342 231024 119398 231033
rect 119342 230959 119398 230968
rect 119356 229094 119384 230959
rect 119080 229066 119384 229094
rect 69478 221776 69534 221785
rect 69478 221711 69534 221720
rect 69386 211576 69442 211585
rect 69386 211511 69442 211520
rect 69400 204950 69428 211511
rect 69388 204944 69440 204950
rect 69388 204886 69440 204892
rect 69294 200696 69350 200705
rect 69294 200631 69350 200640
rect 69308 170406 69336 200631
rect 69388 200388 69440 200394
rect 69388 200330 69440 200336
rect 69400 198150 69428 200330
rect 69388 198144 69440 198150
rect 69388 198086 69440 198092
rect 69492 196654 69520 221711
rect 69662 211984 69718 211993
rect 69662 211919 69718 211928
rect 69572 200048 69624 200054
rect 69572 199990 69624 199996
rect 69584 199646 69612 199990
rect 69572 199640 69624 199646
rect 69572 199582 69624 199588
rect 69480 196648 69532 196654
rect 69480 196590 69532 196596
rect 69676 185638 69704 211919
rect 119080 205634 119108 229066
rect 119342 219600 119398 219609
rect 119342 219535 119398 219544
rect 119160 218476 119212 218482
rect 119160 218418 119212 218424
rect 119172 209774 119200 218418
rect 119356 209774 119384 219535
rect 119448 218006 119476 249630
rect 119724 249150 119752 249750
rect 119712 249144 119764 249150
rect 119712 249086 119764 249092
rect 119712 249008 119764 249014
rect 119712 248950 119764 248956
rect 119724 232762 119752 248950
rect 119712 232756 119764 232762
rect 119712 232698 119764 232704
rect 119816 232558 119844 249766
rect 119908 247722 119936 251767
rect 120000 249014 120028 252554
rect 119988 249008 120040 249014
rect 119988 248950 120040 248956
rect 119896 247716 119948 247722
rect 119896 247658 119948 247664
rect 119804 232552 119856 232558
rect 119804 232494 119856 232500
rect 119896 225004 119948 225010
rect 119896 224946 119948 224952
rect 119528 219428 119580 219434
rect 119528 219370 119580 219376
rect 119540 218521 119568 219370
rect 119526 218512 119582 218521
rect 119526 218447 119528 218456
rect 119580 218447 119582 218456
rect 119528 218418 119580 218424
rect 119436 218000 119488 218006
rect 119436 217942 119488 217948
rect 119172 209746 119292 209774
rect 119356 209746 119476 209774
rect 119080 205606 119200 205634
rect 69768 200382 70058 200410
rect 111260 200394 111288 200763
rect 119172 200530 119200 205606
rect 119160 200524 119212 200530
rect 119160 200466 119212 200472
rect 72608 200388 72660 200394
rect 69768 200190 69796 200382
rect 72608 200330 72660 200336
rect 102830 200388 102882 200394
rect 102830 200330 102882 200336
rect 111248 200388 111300 200394
rect 111248 200330 111300 200336
rect 113180 200388 113232 200394
rect 113180 200330 113232 200336
rect 69848 200320 69900 200326
rect 71274 200320 71326 200326
rect 69848 200262 69900 200268
rect 70674 200288 70730 200297
rect 69756 200184 69808 200190
rect 69756 200126 69808 200132
rect 69860 200114 69888 200262
rect 71274 200262 71326 200268
rect 71286 200237 71314 200262
rect 72620 200237 72648 200330
rect 73252 200320 73304 200326
rect 73252 200262 73304 200268
rect 74540 200320 74592 200326
rect 74540 200262 74592 200268
rect 75184 200320 75236 200326
rect 75184 200262 75236 200268
rect 76472 200320 76524 200326
rect 76472 200262 76524 200268
rect 77116 200320 77168 200326
rect 77116 200262 77168 200268
rect 77760 200320 77812 200326
rect 77760 200262 77812 200268
rect 79048 200320 79100 200326
rect 79048 200262 79100 200268
rect 79692 200320 79744 200326
rect 79692 200262 79744 200268
rect 80980 200320 81032 200326
rect 80980 200262 81032 200268
rect 81624 200320 81676 200326
rect 81624 200262 81676 200268
rect 82912 200320 82964 200326
rect 82912 200262 82964 200268
rect 83556 200320 83608 200326
rect 83556 200262 83608 200268
rect 84200 200320 84252 200326
rect 84200 200262 84252 200268
rect 85488 200320 85540 200326
rect 85488 200262 85540 200268
rect 86132 200320 86184 200326
rect 86132 200262 86184 200268
rect 87420 200320 87472 200326
rect 87420 200262 87472 200268
rect 88064 200320 88116 200326
rect 88064 200262 88116 200268
rect 89352 200320 89404 200326
rect 89352 200262 89404 200268
rect 89996 200320 90048 200326
rect 89996 200262 90048 200268
rect 90640 200320 90692 200326
rect 90640 200262 90692 200268
rect 91928 200320 91980 200326
rect 91928 200262 91980 200268
rect 92572 200320 92624 200326
rect 92572 200262 92624 200268
rect 93860 200320 93912 200326
rect 93860 200262 93912 200268
rect 94504 200320 94556 200326
rect 94504 200262 94556 200268
rect 95792 200320 95844 200326
rect 95792 200262 95844 200268
rect 96436 200320 96488 200326
rect 96436 200262 96488 200268
rect 97724 200320 97776 200326
rect 97724 200262 97776 200268
rect 98368 200320 98420 200326
rect 98368 200262 98420 200268
rect 99012 200320 99064 200326
rect 99012 200262 99064 200268
rect 100300 200320 100352 200326
rect 100300 200262 100352 200268
rect 100898 200320 100950 200326
rect 100898 200262 100950 200268
rect 102232 200320 102284 200326
rect 102232 200262 102284 200268
rect 73264 200237 73292 200262
rect 74552 200237 74580 200262
rect 75196 200237 75224 200262
rect 76484 200237 76512 200262
rect 77128 200237 77156 200262
rect 77772 200237 77800 200262
rect 79060 200237 79088 200262
rect 79704 200237 79732 200262
rect 80992 200237 81020 200262
rect 81636 200237 81664 200262
rect 82924 200237 82952 200262
rect 83568 200237 83596 200262
rect 84212 200237 84240 200262
rect 85500 200237 85528 200262
rect 86144 200237 86172 200262
rect 87432 200237 87460 200262
rect 88076 200237 88104 200262
rect 89364 200237 89392 200262
rect 90008 200237 90036 200262
rect 90652 200237 90680 200262
rect 91940 200237 91968 200262
rect 92584 200237 92612 200262
rect 93872 200237 93900 200262
rect 94516 200237 94544 200262
rect 95804 200237 95832 200262
rect 96448 200237 96476 200262
rect 97736 200237 97764 200262
rect 98380 200237 98408 200262
rect 99024 200237 99052 200262
rect 100312 200237 100340 200262
rect 100910 200237 100938 200262
rect 102244 200237 102272 200262
rect 102842 200237 102870 200330
rect 104164 200320 104216 200326
rect 104164 200262 104216 200268
rect 104808 200320 104860 200326
rect 104808 200262 104860 200268
rect 105406 200320 105458 200326
rect 105406 200262 105458 200268
rect 106740 200320 106792 200326
rect 106740 200262 106792 200268
rect 107384 200320 107436 200326
rect 107384 200262 107436 200268
rect 108672 200320 108724 200326
rect 108672 200262 108724 200268
rect 109316 200320 109368 200326
rect 109316 200262 109368 200268
rect 110604 200320 110656 200326
rect 110604 200262 110656 200268
rect 111892 200320 111944 200326
rect 111892 200262 111944 200268
rect 104176 200237 104204 200262
rect 104820 200237 104848 200262
rect 105418 200237 105446 200262
rect 106752 200237 106780 200262
rect 107396 200237 107424 200262
rect 108684 200237 108712 200262
rect 109328 200237 109356 200262
rect 110616 200237 110644 200262
rect 111904 200237 111932 200262
rect 113192 200237 113220 200330
rect 113778 200320 113830 200326
rect 113778 200262 113830 200268
rect 115112 200320 115164 200326
rect 115112 200262 115164 200268
rect 115756 200320 115808 200326
rect 115756 200262 115808 200268
rect 117044 200320 117096 200326
rect 117044 200262 117096 200268
rect 117688 200320 117740 200326
rect 117688 200262 117740 200268
rect 113790 200237 113818 200262
rect 115124 200237 115152 200262
rect 115768 200237 115796 200262
rect 117056 200237 117084 200262
rect 117700 200237 117728 200262
rect 119002 200246 119200 200274
rect 70674 200223 70730 200232
rect 119068 200116 119120 200122
rect 69860 200086 69980 200114
rect 69952 200002 69980 200086
rect 119068 200058 119120 200064
rect 69952 199974 70440 200002
rect 70308 196648 70360 196654
rect 70308 196590 70360 196596
rect 69664 185632 69716 185638
rect 69664 185574 69716 185580
rect 69388 175976 69440 175982
rect 69386 175944 69388 175953
rect 69440 175944 69442 175953
rect 69386 175879 69442 175888
rect 69296 170400 69348 170406
rect 69296 170342 69348 170348
rect 69572 115048 69624 115054
rect 69572 114990 69624 114996
rect 69388 113824 69440 113830
rect 69388 113766 69440 113772
rect 69400 113422 69428 113766
rect 69388 113416 69440 113422
rect 69388 113358 69440 113364
rect 69296 111784 69348 111790
rect 69296 111726 69348 111732
rect 69204 111716 69256 111722
rect 69204 111658 69256 111664
rect 69110 106040 69166 106049
rect 69110 105975 69166 105984
rect 69018 89040 69074 89049
rect 69018 88975 69074 88984
rect 68834 86320 68890 86329
rect 68834 86255 68890 86264
rect 68848 74534 68876 86255
rect 68926 75848 68982 75857
rect 68926 75783 68982 75792
rect 68940 74905 68968 75783
rect 68926 74896 68982 74905
rect 68926 74831 68982 74840
rect 68756 74506 68876 74534
rect 68650 71360 68706 71369
rect 68650 71295 68706 71304
rect 68560 69760 68612 69766
rect 68560 69702 68612 69708
rect 68466 67280 68522 67289
rect 68466 67215 68522 67224
rect 68282 65784 68338 65793
rect 68282 65719 68338 65728
rect 68756 65414 68784 74506
rect 68834 74080 68890 74089
rect 68834 74015 68890 74024
rect 68848 67386 68876 74015
rect 68836 67380 68888 67386
rect 68836 67322 68888 67328
rect 68940 66706 68968 74831
rect 68928 66700 68980 66706
rect 68928 66642 68980 66648
rect 68744 65408 68796 65414
rect 68744 65350 68796 65356
rect 67548 64728 67600 64734
rect 67548 64670 67600 64676
rect 65524 33108 65576 33114
rect 65524 33050 65576 33056
rect 3516 20664 3568 20670
rect 3516 20606 3568 20612
rect 3528 19417 3556 20606
rect 3514 19408 3570 19417
rect 3514 19343 3570 19352
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4172 2854 4200 4762
rect 69124 3466 69152 105975
rect 69204 96552 69256 96558
rect 69204 96494 69256 96500
rect 69216 95305 69244 96494
rect 69202 95296 69258 95305
rect 69202 95231 69258 95240
rect 69216 69737 69244 95231
rect 69308 87009 69336 111726
rect 69400 90545 69428 113358
rect 69480 112532 69532 112538
rect 69480 112474 69532 112480
rect 69492 93945 69520 112474
rect 69584 99385 69612 114990
rect 70216 114708 70268 114714
rect 70216 114650 70268 114656
rect 69664 112260 69716 112266
rect 69664 112202 69716 112208
rect 69570 99376 69626 99385
rect 69570 99311 69626 99320
rect 69676 97345 69704 112202
rect 70032 111988 70084 111994
rect 70032 111930 70084 111936
rect 70044 111724 70072 111930
rect 69848 111716 69900 111722
rect 69848 111658 69900 111664
rect 69860 111625 69888 111658
rect 69846 111616 69902 111625
rect 69846 111551 69902 111560
rect 70228 108633 70256 114650
rect 70320 113626 70348 196590
rect 70308 113620 70360 113626
rect 70308 113562 70360 113568
rect 70320 111790 70348 113562
rect 70308 111784 70360 111790
rect 70308 111726 70360 111732
rect 70308 110492 70360 110498
rect 70308 110434 70360 110440
rect 70320 109993 70348 110434
rect 70306 109984 70362 109993
rect 70306 109919 70362 109928
rect 70214 108624 70270 108633
rect 70214 108559 70270 108568
rect 69662 97336 69718 97345
rect 69662 97271 69718 97280
rect 69478 93936 69534 93945
rect 69478 93871 69534 93880
rect 69386 90536 69442 90545
rect 69386 90471 69442 90480
rect 69294 87000 69350 87009
rect 69294 86935 69350 86944
rect 69294 82240 69350 82249
rect 69294 82175 69350 82184
rect 69202 69728 69258 69737
rect 69202 69663 69258 69672
rect 69308 65482 69336 82175
rect 69754 80200 69810 80209
rect 69754 80135 69810 80144
rect 69386 79520 69442 79529
rect 69386 79455 69442 79464
rect 69296 65476 69348 65482
rect 69296 65418 69348 65424
rect 69400 64258 69428 79455
rect 69478 76800 69534 76809
rect 69478 76735 69534 76744
rect 69492 64666 69520 76735
rect 69570 73264 69626 73273
rect 69570 73199 69626 73208
rect 69584 72729 69612 73199
rect 69570 72720 69626 72729
rect 69570 72655 69626 72664
rect 69584 64841 69612 72655
rect 69662 70680 69718 70689
rect 69662 70615 69718 70624
rect 69570 64832 69626 64841
rect 69570 64767 69626 64776
rect 69480 64660 69532 64666
rect 69480 64602 69532 64608
rect 69676 64530 69704 70615
rect 69768 64598 69796 80135
rect 69846 71360 69902 71369
rect 69846 71295 69902 71304
rect 69756 64592 69808 64598
rect 69756 64534 69808 64540
rect 69664 64524 69716 64530
rect 69664 64466 69716 64472
rect 69860 64394 69888 71295
rect 70412 70310 70440 199974
rect 73160 199980 73212 199986
rect 73160 199922 73212 199928
rect 73252 199980 73304 199986
rect 73252 199922 73304 199928
rect 74540 199980 74592 199986
rect 74540 199922 74592 199928
rect 75092 199980 75144 199986
rect 75092 199922 75144 199928
rect 76472 199980 76524 199986
rect 76472 199922 76524 199928
rect 77116 199980 77168 199986
rect 77116 199922 77168 199928
rect 77760 199980 77812 199986
rect 77760 199922 77812 199928
rect 79048 199980 79100 199986
rect 79048 199922 79100 199928
rect 79692 199980 79744 199986
rect 79692 199922 79744 199928
rect 80980 199980 81032 199986
rect 80980 199922 81032 199928
rect 81624 199980 81676 199986
rect 81624 199922 81676 199928
rect 82912 199980 82964 199986
rect 82912 199922 82964 199928
rect 83556 199980 83608 199986
rect 83556 199922 83608 199928
rect 84200 199980 84252 199986
rect 84200 199922 84252 199928
rect 85488 199980 85540 199986
rect 85488 199922 85540 199928
rect 86132 199980 86184 199986
rect 86132 199922 86184 199928
rect 87420 199980 87472 199986
rect 87420 199922 87472 199928
rect 87972 199980 88024 199986
rect 87972 199922 88024 199928
rect 89352 199980 89404 199986
rect 89352 199922 89404 199928
rect 89904 199980 89956 199986
rect 89904 199922 89956 199928
rect 90640 199980 90692 199986
rect 90640 199922 90692 199928
rect 91836 199980 91888 199986
rect 91836 199922 91888 199928
rect 92480 199980 92532 199986
rect 92480 199922 92532 199928
rect 93860 199980 93912 199986
rect 93860 199922 93912 199928
rect 94412 199980 94464 199986
rect 94412 199922 94464 199928
rect 95700 199980 95752 199986
rect 95700 199922 95752 199928
rect 96436 199980 96488 199986
rect 96436 199922 96488 199928
rect 97264 199980 97316 199986
rect 97264 199922 97316 199928
rect 98276 199980 98328 199986
rect 98276 199922 98328 199928
rect 98552 199980 98604 199986
rect 98552 199922 98604 199928
rect 98920 199980 98972 199986
rect 98920 199922 98972 199928
rect 100300 199980 100352 199986
rect 100300 199922 100352 199928
rect 101312 199980 101364 199986
rect 101312 199922 101364 199928
rect 103428 199980 103480 199986
rect 103428 199922 103480 199928
rect 104164 199980 104216 199986
rect 104164 199922 104216 199928
rect 104256 199980 104308 199986
rect 104256 199922 104308 199928
rect 104808 199980 104860 199986
rect 104808 199922 104860 199928
rect 105360 199980 105412 199986
rect 105360 199922 105412 199928
rect 107476 199980 107528 199986
rect 107476 199922 107528 199928
rect 108764 199980 108816 199986
rect 108764 199922 108816 199928
rect 109316 199980 109368 199986
rect 109316 199922 109368 199928
rect 111248 199980 111300 199986
rect 111248 199922 111300 199928
rect 112536 199980 112588 199986
rect 112536 199922 112588 199928
rect 113180 199980 113232 199986
rect 113180 199922 113232 199928
rect 114468 199980 114520 199986
rect 114468 199922 114520 199928
rect 115296 199980 115348 199986
rect 115296 199922 115348 199928
rect 115848 199980 115900 199986
rect 115848 199922 115900 199928
rect 116584 199980 116636 199986
rect 116584 199922 116636 199928
rect 117320 199980 117372 199986
rect 117320 199922 117372 199928
rect 117688 199980 117740 199986
rect 117688 199922 117740 199928
rect 70490 199880 70546 199889
rect 70490 199815 70546 199824
rect 70504 171834 70532 199815
rect 73172 199374 73200 199922
rect 72700 199368 72752 199374
rect 72700 199310 72752 199316
rect 73160 199368 73212 199374
rect 73160 199310 73212 199316
rect 72606 198792 72662 198801
rect 71044 198756 71096 198762
rect 72606 198727 72662 198736
rect 71044 198698 71096 198704
rect 71056 180130 71084 198698
rect 72620 183530 72648 198727
rect 72712 186998 72740 199310
rect 72700 186992 72752 186998
rect 72700 186934 72752 186940
rect 72608 183524 72660 183530
rect 72608 183466 72660 183472
rect 71044 180124 71096 180130
rect 71044 180066 71096 180072
rect 70492 171828 70544 171834
rect 70492 171770 70544 171776
rect 70504 70666 70532 171770
rect 73264 169386 73292 199922
rect 73252 169380 73304 169386
rect 73252 169322 73304 169328
rect 74552 169017 74580 199922
rect 74828 199714 75040 199730
rect 74816 199708 75052 199714
rect 74868 199702 75000 199708
rect 74816 199650 74868 199656
rect 75000 199650 75052 199656
rect 74724 199640 74776 199646
rect 74724 199582 74776 199588
rect 74736 199238 74764 199582
rect 74724 199232 74776 199238
rect 74724 199174 74776 199180
rect 75104 198422 75132 199922
rect 75184 199912 75236 199918
rect 75184 199854 75236 199860
rect 75196 199306 75224 199854
rect 75276 199776 75328 199782
rect 75276 199718 75328 199724
rect 75288 199646 75316 199718
rect 75276 199640 75328 199646
rect 75276 199582 75328 199588
rect 75184 199300 75236 199306
rect 75184 199242 75236 199248
rect 75092 198416 75144 198422
rect 75092 198358 75144 198364
rect 75104 195974 75132 198358
rect 76484 196790 76512 199922
rect 77128 197878 77156 199922
rect 77116 197872 77168 197878
rect 77116 197814 77168 197820
rect 76472 196784 76524 196790
rect 76472 196726 76524 196732
rect 75104 195946 75224 195974
rect 75196 170474 75224 195946
rect 77772 181490 77800 199922
rect 79060 198218 79088 199922
rect 79048 198212 79100 198218
rect 79048 198154 79100 198160
rect 79704 198082 79732 199922
rect 79692 198076 79744 198082
rect 79692 198018 79744 198024
rect 79324 197872 79376 197878
rect 79324 197814 79376 197820
rect 77760 181484 77812 181490
rect 77760 181426 77812 181432
rect 75184 170468 75236 170474
rect 75184 170410 75236 170416
rect 79336 169318 79364 197814
rect 80992 173262 81020 199922
rect 81636 198422 81664 199922
rect 82082 199336 82138 199345
rect 82082 199271 82084 199280
rect 82136 199271 82138 199280
rect 82084 199242 82136 199248
rect 81624 198416 81676 198422
rect 81624 198358 81676 198364
rect 82924 184210 82952 199922
rect 82912 184204 82964 184210
rect 82912 184146 82964 184152
rect 80980 173256 81032 173262
rect 80980 173198 81032 173204
rect 83568 170610 83596 199922
rect 83556 170604 83608 170610
rect 83556 170546 83608 170552
rect 79324 169312 79376 169318
rect 79324 169254 79376 169260
rect 84212 169114 84240 199922
rect 84660 199912 84712 199918
rect 84660 199854 84712 199860
rect 84672 199238 84700 199854
rect 84844 199844 84896 199850
rect 84844 199786 84896 199792
rect 84752 199368 84804 199374
rect 84752 199310 84804 199316
rect 84764 199238 84792 199310
rect 84660 199232 84712 199238
rect 84660 199174 84712 199180
rect 84752 199232 84804 199238
rect 84752 199174 84804 199180
rect 84856 199170 84884 199786
rect 84936 199368 84988 199374
rect 84934 199336 84936 199345
rect 84988 199336 84990 199345
rect 84934 199271 84990 199280
rect 84844 199164 84896 199170
rect 84844 199106 84896 199112
rect 85500 198082 85528 199922
rect 85488 198076 85540 198082
rect 85488 198018 85540 198024
rect 86144 197946 86172 199922
rect 87432 198626 87460 199922
rect 87420 198620 87472 198626
rect 87420 198562 87472 198568
rect 86132 197940 86184 197946
rect 86132 197882 86184 197888
rect 86224 196784 86276 196790
rect 86224 196726 86276 196732
rect 84200 169108 84252 169114
rect 84200 169050 84252 169056
rect 74538 169008 74594 169017
rect 74538 168943 74594 168952
rect 86236 167686 86264 196726
rect 87432 195974 87460 198562
rect 87432 195946 87644 195974
rect 87616 169182 87644 195946
rect 87984 195294 88012 199922
rect 87972 195288 88024 195294
rect 87972 195230 88024 195236
rect 89364 189854 89392 199922
rect 89916 197878 89944 199922
rect 89904 197872 89956 197878
rect 89904 197814 89956 197820
rect 89352 189848 89404 189854
rect 89352 189790 89404 189796
rect 90652 182850 90680 199922
rect 91848 198626 91876 199922
rect 91836 198620 91888 198626
rect 91836 198562 91888 198568
rect 92492 197402 92520 199922
rect 93872 198121 93900 199922
rect 93858 198112 93914 198121
rect 93858 198047 93914 198056
rect 92480 197396 92532 197402
rect 92480 197338 92532 197344
rect 94424 195362 94452 199922
rect 95712 198218 95740 199922
rect 95700 198212 95752 198218
rect 95700 198154 95752 198160
rect 94596 197396 94648 197402
rect 94596 197338 94648 197344
rect 94412 195356 94464 195362
rect 94412 195298 94464 195304
rect 90640 182844 90692 182850
rect 90640 182786 90692 182792
rect 94608 169250 94636 197338
rect 96448 170678 96476 199922
rect 97276 198490 97304 199922
rect 97264 198484 97316 198490
rect 97264 198426 97316 198432
rect 97276 177410 97304 198426
rect 98288 195430 98316 199922
rect 98564 199306 98592 199922
rect 98644 199844 98696 199850
rect 98644 199786 98696 199792
rect 98552 199300 98604 199306
rect 98552 199242 98604 199248
rect 98656 199238 98684 199786
rect 98736 199776 98788 199782
rect 98736 199718 98788 199724
rect 98748 199374 98776 199718
rect 98736 199368 98788 199374
rect 98736 199310 98788 199316
rect 98644 199232 98696 199238
rect 98644 199174 98696 199180
rect 98932 198490 98960 199922
rect 98920 198484 98972 198490
rect 98920 198426 98972 198432
rect 100312 195498 100340 199922
rect 101324 198354 101352 199922
rect 103440 198529 103468 199922
rect 104072 198552 104124 198558
rect 103426 198520 103482 198529
rect 104072 198494 104124 198500
rect 103426 198455 103482 198464
rect 101312 198348 101364 198354
rect 101312 198290 101364 198296
rect 100300 195492 100352 195498
rect 100300 195434 100352 195440
rect 98276 195424 98328 195430
rect 98276 195366 98328 195372
rect 97264 177404 97316 177410
rect 97264 177346 97316 177352
rect 96436 170672 96488 170678
rect 96436 170614 96488 170620
rect 94596 169244 94648 169250
rect 94596 169186 94648 169192
rect 87604 169176 87656 169182
rect 87604 169118 87656 169124
rect 103440 169046 103468 198455
rect 104084 197810 104112 198494
rect 104072 197804 104124 197810
rect 104072 197746 104124 197752
rect 104176 197674 104204 199922
rect 104268 198286 104296 199922
rect 104256 198280 104308 198286
rect 104256 198222 104308 198228
rect 104820 197742 104848 199922
rect 104808 197736 104860 197742
rect 104808 197678 104860 197684
rect 104164 197668 104216 197674
rect 104164 197610 104216 197616
rect 105372 195566 105400 199922
rect 107200 199844 107252 199850
rect 107200 199786 107252 199792
rect 106280 198484 106332 198490
rect 106280 198426 106332 198432
rect 105360 195560 105412 195566
rect 105360 195502 105412 195508
rect 103428 169040 103480 169046
rect 103428 168982 103480 168988
rect 86224 167680 86276 167686
rect 86224 167622 86276 167628
rect 95884 123480 95936 123486
rect 95884 123422 95936 123428
rect 88340 122460 88392 122466
rect 88340 122402 88392 122408
rect 83096 121168 83148 121174
rect 83096 121110 83148 121116
rect 80520 120964 80572 120970
rect 80520 120906 80572 120912
rect 79324 119536 79376 119542
rect 79324 119478 79376 119484
rect 78496 119468 78548 119474
rect 78496 119410 78548 119416
rect 78508 118658 78536 119410
rect 78588 119400 78640 119406
rect 78588 119342 78640 119348
rect 78496 118652 78548 118658
rect 78496 118594 78548 118600
rect 77760 118584 77812 118590
rect 77760 118526 77812 118532
rect 76470 118008 76526 118017
rect 76470 117943 76526 117952
rect 75920 117428 75972 117434
rect 75920 117370 75972 117376
rect 75932 117230 75960 117370
rect 76484 117298 76512 117943
rect 76472 117292 76524 117298
rect 76472 117234 76524 117240
rect 77116 117292 77168 117298
rect 77116 117234 77168 117240
rect 75920 117224 75972 117230
rect 75920 117166 75972 117172
rect 73250 116240 73306 116249
rect 73250 116175 73306 116184
rect 72608 116136 72660 116142
rect 72608 116078 72660 116084
rect 71688 114912 71740 114918
rect 71688 114854 71740 114860
rect 71700 114374 71728 114854
rect 71320 114368 71372 114374
rect 71320 114310 71372 114316
rect 71688 114368 71740 114374
rect 71688 114310 71740 114316
rect 70676 111920 70728 111926
rect 70676 111862 70728 111868
rect 70688 111724 70716 111862
rect 71332 111724 71360 114310
rect 71964 114232 72016 114238
rect 71964 114174 72016 114180
rect 71596 112464 71648 112470
rect 71596 112406 71648 112412
rect 71608 111926 71636 112406
rect 71596 111920 71648 111926
rect 71596 111862 71648 111868
rect 71976 111724 72004 114174
rect 72332 113620 72384 113626
rect 72332 113562 72384 113568
rect 72344 113490 72372 113562
rect 72332 113484 72384 113490
rect 72332 113426 72384 113432
rect 72620 111724 72648 116078
rect 73068 114980 73120 114986
rect 73068 114922 73120 114928
rect 73080 114238 73108 114922
rect 73068 114232 73120 114238
rect 73068 114174 73120 114180
rect 73264 111724 73292 116175
rect 75552 115320 75604 115326
rect 75552 115262 75604 115268
rect 74540 114368 74592 114374
rect 74540 114310 74592 114316
rect 74552 111724 74580 114310
rect 74998 112160 75054 112169
rect 74998 112095 75054 112104
rect 75012 111897 75040 112095
rect 75184 112056 75236 112062
rect 75236 112004 75316 112010
rect 75184 111998 75316 112004
rect 75196 111982 75316 111998
rect 74998 111888 75054 111897
rect 75288 111874 75316 111982
rect 75460 111920 75512 111926
rect 75288 111868 75460 111874
rect 75288 111862 75512 111868
rect 75288 111846 75500 111862
rect 74998 111823 75054 111832
rect 75564 111738 75592 115262
rect 75828 115252 75880 115258
rect 75828 115194 75880 115200
rect 75840 114442 75868 115194
rect 75828 114436 75880 114442
rect 75828 114378 75880 114384
rect 75644 112056 75696 112062
rect 75644 111998 75696 112004
rect 75210 111710 75592 111738
rect 75656 111722 75684 111998
rect 75840 111724 75868 114378
rect 75932 114374 75960 117166
rect 76470 116512 76526 116521
rect 76470 116447 76526 116456
rect 75920 114368 75972 114374
rect 75920 114310 75972 114316
rect 76484 111724 76512 116447
rect 77128 111724 77156 117234
rect 77772 111724 77800 118526
rect 78508 111738 78536 118594
rect 78600 118590 78628 119342
rect 78588 118584 78640 118590
rect 78588 118526 78640 118532
rect 79336 114510 79364 119478
rect 80060 117496 80112 117502
rect 80060 117438 80112 117444
rect 80072 115326 80100 117438
rect 80060 115320 80112 115326
rect 80060 115262 80112 115268
rect 79324 114504 79376 114510
rect 79324 114446 79376 114452
rect 79336 111738 79364 114446
rect 79692 113688 79744 113694
rect 79692 113630 79744 113636
rect 75644 111716 75696 111722
rect 78430 111710 78536 111738
rect 79074 111710 79364 111738
rect 79704 111724 79732 113630
rect 80532 111738 80560 120906
rect 82912 116612 82964 116618
rect 82912 116554 82964 116560
rect 82268 115320 82320 115326
rect 82268 115262 82320 115268
rect 81624 113960 81676 113966
rect 81624 113902 81676 113908
rect 80532 111710 81006 111738
rect 81636 111724 81664 113902
rect 82280 111724 82308 115262
rect 82924 111724 82952 116554
rect 83108 111738 83136 121110
rect 85580 121100 85632 121106
rect 85580 121042 85632 121048
rect 84200 120828 84252 120834
rect 84200 120770 84252 120776
rect 83108 111710 83582 111738
rect 84212 111724 84240 120770
rect 84384 116680 84436 116686
rect 84384 116622 84436 116628
rect 84396 111738 84424 116622
rect 85592 113174 85620 121042
rect 86868 120760 86920 120766
rect 86868 120702 86920 120708
rect 86132 114096 86184 114102
rect 86132 114038 86184 114044
rect 85500 113146 85620 113174
rect 84396 111710 84870 111738
rect 85500 111724 85528 113146
rect 86144 111724 86172 114038
rect 86880 113694 86908 120702
rect 86960 119672 87012 119678
rect 86960 119614 87012 119620
rect 86868 113688 86920 113694
rect 86868 113630 86920 113636
rect 86972 111738 87000 119614
rect 88352 113174 88380 122402
rect 92204 122392 92256 122398
rect 92204 122334 92256 122340
rect 91100 122188 91152 122194
rect 91100 122130 91152 122136
rect 89720 119604 89772 119610
rect 89720 119546 89772 119552
rect 88708 113892 88760 113898
rect 88708 113834 88760 113840
rect 88260 113146 88380 113174
rect 88260 111738 88288 113146
rect 86972 111710 87446 111738
rect 88090 111710 88288 111738
rect 88720 111724 88748 113834
rect 89352 113824 89404 113830
rect 89352 113766 89404 113772
rect 89364 111724 89392 113766
rect 89732 111738 89760 119546
rect 90640 114436 90692 114442
rect 90640 114378 90692 114384
rect 89732 111710 90022 111738
rect 90652 111724 90680 114378
rect 91112 111738 91140 122130
rect 91560 118040 91612 118046
rect 91560 117982 91612 117988
rect 91572 111738 91600 117982
rect 92216 114442 92244 122334
rect 93860 122256 93912 122262
rect 93860 122198 93912 122204
rect 92480 118108 92532 118114
rect 92480 118050 92532 118056
rect 92204 114436 92256 114442
rect 92204 114378 92256 114384
rect 92492 113174 92520 118050
rect 92492 113146 92612 113174
rect 91112 111710 91310 111738
rect 91572 111710 91954 111738
rect 92584 111724 92612 113146
rect 93872 111724 93900 122198
rect 95424 121304 95476 121310
rect 95424 121246 95476 121252
rect 94136 121032 94188 121038
rect 94136 120974 94188 120980
rect 94148 111738 94176 120974
rect 95148 114164 95200 114170
rect 95148 114106 95200 114112
rect 94148 111710 94530 111738
rect 95160 111724 95188 114106
rect 95436 111738 95464 121246
rect 95896 114510 95924 123422
rect 99288 122324 99340 122330
rect 99288 122266 99340 122272
rect 98000 116748 98052 116754
rect 98000 116690 98052 116696
rect 97724 115932 97776 115938
rect 97724 115874 97776 115880
rect 97080 115388 97132 115394
rect 97080 115330 97132 115336
rect 95884 114504 95936 114510
rect 95884 114446 95936 114452
rect 96436 114504 96488 114510
rect 96436 114446 96488 114452
rect 95436 111710 95818 111738
rect 96448 111724 96476 114446
rect 97092 111724 97120 115330
rect 97736 111724 97764 115874
rect 98012 111738 98040 116690
rect 99300 115938 99328 122266
rect 104900 121644 104952 121650
rect 104900 121586 104952 121592
rect 102416 121440 102468 121446
rect 102416 121382 102468 121388
rect 102140 121236 102192 121242
rect 102140 121178 102192 121184
rect 99840 117972 99892 117978
rect 99840 117914 99892 117920
rect 99288 115932 99340 115938
rect 99288 115874 99340 115880
rect 99012 114028 99064 114034
rect 99012 113970 99064 113976
rect 98012 111710 98394 111738
rect 99024 111724 99052 113970
rect 99852 111738 99880 117914
rect 100944 114300 100996 114306
rect 100944 114242 100996 114248
rect 100760 111852 100812 111858
rect 100760 111794 100812 111800
rect 100772 111738 100800 111794
rect 100956 111738 100984 114242
rect 101588 114232 101640 114238
rect 101588 114174 101640 114180
rect 101600 111926 101628 114174
rect 102152 113174 102180 121178
rect 102152 113146 102272 113174
rect 101588 111920 101640 111926
rect 101588 111862 101640 111868
rect 99852 111710 100326 111738
rect 100772 111724 100984 111738
rect 101600 111724 101628 111862
rect 102244 111724 102272 113146
rect 102428 111738 102456 121382
rect 103796 121372 103848 121378
rect 103796 121314 103848 121320
rect 103612 119740 103664 119746
rect 103612 119682 103664 119688
rect 103624 111738 103652 119682
rect 100772 111710 100970 111724
rect 102428 111710 102902 111738
rect 103546 111710 103652 111738
rect 103808 111738 103836 121314
rect 104912 115818 104940 121586
rect 104820 115790 104940 115818
rect 103808 111710 104190 111738
rect 104820 111724 104848 115790
rect 105478 111722 105768 111738
rect 105478 111716 105780 111722
rect 105478 111710 105728 111716
rect 75644 111658 75696 111664
rect 105728 111658 105780 111664
rect 106186 77208 106242 77217
rect 106186 77143 106242 77152
rect 106200 76537 106228 77143
rect 106186 76528 106242 76537
rect 106186 76463 106242 76472
rect 106186 75032 106242 75041
rect 106016 74990 106186 75018
rect 106016 71754 106044 74990
rect 106186 74967 106242 74976
rect 106188 74588 106240 74594
rect 106188 74530 106240 74536
rect 106096 73228 106148 73234
rect 106096 73170 106148 73176
rect 106108 71874 106136 73170
rect 106200 71874 106228 74530
rect 106096 71868 106148 71874
rect 106096 71810 106148 71816
rect 106188 71868 106240 71874
rect 106188 71810 106240 71816
rect 106016 71726 106228 71754
rect 106096 71596 106148 71602
rect 106096 71538 106148 71544
rect 106004 70780 106056 70786
rect 106004 70722 106056 70728
rect 70504 70638 70702 70666
rect 70400 70304 70452 70310
rect 70400 70246 70452 70252
rect 70044 70106 70072 70244
rect 70032 70100 70084 70106
rect 70032 70042 70084 70048
rect 70306 70000 70362 70009
rect 70306 69935 70362 69944
rect 70320 69834 70348 69935
rect 70308 69828 70360 69834
rect 70308 69770 70360 69776
rect 70412 67969 70440 70246
rect 70504 68066 70532 70638
rect 74540 70440 74592 70446
rect 74540 70382 74592 70388
rect 75184 70440 75236 70446
rect 75184 70382 75236 70388
rect 76472 70440 76524 70446
rect 76472 70382 76524 70388
rect 71274 70304 71326 70310
rect 71274 70246 71326 70252
rect 71964 70304 72016 70310
rect 71964 70246 72016 70252
rect 72608 70304 72660 70310
rect 72608 70246 72660 70252
rect 73252 70304 73304 70310
rect 73252 70246 73304 70252
rect 73896 70304 73948 70310
rect 73896 70246 73948 70252
rect 71286 70244 71314 70246
rect 71976 70244 72004 70246
rect 72620 70244 72648 70246
rect 73264 70244 73292 70246
rect 73908 70244 73936 70246
rect 74552 70244 74580 70382
rect 75196 70244 75224 70382
rect 76484 70244 76512 70382
rect 82872 70372 82924 70378
rect 82872 70314 82924 70320
rect 100944 70372 100996 70378
rect 100944 70314 100996 70320
rect 77116 70304 77168 70310
rect 77116 70246 77168 70252
rect 77760 70304 77812 70310
rect 77760 70246 77812 70252
rect 78404 70304 78456 70310
rect 78404 70246 78456 70252
rect 79048 70304 79100 70310
rect 79048 70246 79100 70252
rect 79692 70304 79744 70310
rect 79692 70246 79744 70252
rect 80336 70304 80388 70310
rect 80336 70246 80388 70252
rect 80980 70304 81032 70310
rect 80980 70246 81032 70252
rect 81624 70304 81676 70310
rect 81624 70246 81676 70252
rect 77128 70244 77156 70246
rect 77772 70244 77800 70246
rect 78416 70244 78444 70246
rect 79060 70244 79088 70246
rect 79704 70244 79732 70246
rect 80348 70244 80376 70246
rect 80992 70244 81020 70246
rect 81636 70244 81664 70246
rect 82884 70244 82912 70314
rect 83556 70304 83608 70310
rect 83556 70246 83608 70252
rect 84200 70304 84252 70310
rect 84200 70246 84252 70252
rect 84860 70304 84912 70310
rect 84860 70246 84912 70252
rect 85488 70304 85540 70310
rect 85488 70246 85540 70252
rect 86132 70304 86184 70310
rect 86132 70246 86184 70252
rect 86776 70304 86828 70310
rect 86776 70246 86828 70252
rect 87420 70304 87472 70310
rect 87420 70246 87472 70252
rect 88064 70304 88116 70310
rect 88064 70246 88116 70252
rect 89352 70304 89404 70310
rect 89352 70246 89404 70252
rect 89996 70304 90048 70310
rect 89996 70246 90048 70252
rect 90640 70304 90692 70310
rect 90640 70246 90692 70252
rect 91284 70304 91336 70310
rect 91284 70246 91336 70252
rect 91928 70304 91980 70310
rect 91928 70246 91980 70252
rect 92572 70304 92624 70310
rect 92572 70246 92624 70252
rect 93216 70304 93268 70310
rect 93216 70246 93268 70252
rect 93860 70304 93912 70310
rect 93860 70246 93912 70252
rect 94520 70304 94572 70310
rect 94520 70246 94572 70252
rect 95792 70304 95844 70310
rect 95792 70246 95844 70252
rect 96436 70304 96488 70310
rect 96436 70246 96488 70252
rect 97080 70304 97132 70310
rect 97080 70246 97132 70252
rect 97724 70304 97776 70310
rect 97724 70246 97776 70252
rect 98368 70304 98420 70310
rect 98368 70246 98420 70252
rect 99012 70304 99064 70310
rect 99012 70246 99064 70252
rect 99656 70304 99708 70310
rect 99656 70246 99708 70252
rect 100300 70304 100352 70310
rect 100300 70246 100352 70252
rect 83568 70244 83596 70246
rect 84212 70244 84240 70246
rect 84872 70244 84900 70246
rect 85500 70244 85528 70246
rect 86144 70244 86172 70246
rect 86788 70244 86816 70246
rect 87432 70244 87460 70246
rect 88076 70244 88104 70246
rect 89364 70244 89392 70246
rect 90008 70244 90036 70246
rect 90652 70244 90680 70246
rect 91296 70244 91324 70246
rect 91940 70244 91968 70246
rect 92584 70244 92612 70246
rect 93228 70244 93256 70246
rect 93872 70244 93900 70246
rect 94532 70244 94560 70246
rect 95804 70244 95832 70246
rect 96448 70244 96476 70246
rect 97092 70244 97120 70246
rect 97736 70244 97764 70246
rect 98380 70244 98408 70246
rect 99024 70244 99052 70246
rect 99668 70244 99696 70246
rect 100312 70244 100340 70246
rect 100956 70244 100984 70314
rect 102232 70304 102284 70310
rect 102232 70246 102284 70252
rect 102876 70304 102928 70310
rect 102876 70246 102928 70252
rect 103520 70304 103572 70310
rect 103520 70246 103572 70252
rect 104180 70304 104232 70310
rect 104180 70246 104232 70252
rect 104824 70304 104876 70310
rect 104824 70246 104876 70252
rect 105468 70304 105520 70310
rect 105468 70246 105520 70252
rect 102244 70244 102272 70246
rect 102888 70244 102916 70246
rect 103532 70244 103560 70246
rect 104192 70244 104220 70246
rect 104836 70244 104864 70246
rect 105480 70244 105508 70246
rect 71964 69964 72016 69970
rect 71964 69906 72016 69912
rect 72608 69964 72660 69970
rect 72608 69906 72660 69912
rect 73344 69964 73396 69970
rect 73344 69906 73396 69912
rect 73988 69964 74040 69970
rect 73988 69906 74040 69912
rect 74540 69964 74592 69970
rect 74540 69906 74592 69912
rect 75184 69964 75236 69970
rect 75184 69906 75236 69912
rect 76564 69964 76616 69970
rect 76564 69906 76616 69912
rect 77116 69964 77168 69970
rect 77116 69906 77168 69912
rect 77760 69964 77812 69970
rect 77760 69906 77812 69912
rect 78404 69964 78456 69970
rect 78404 69906 78456 69912
rect 79048 69964 79100 69970
rect 79048 69906 79100 69912
rect 79692 69964 79744 69970
rect 79692 69906 79744 69912
rect 80428 69964 80480 69970
rect 80428 69906 80480 69912
rect 81072 69964 81124 69970
rect 81072 69906 81124 69912
rect 81716 69964 81768 69970
rect 81716 69906 81768 69912
rect 82912 69964 82964 69970
rect 82912 69906 82964 69912
rect 83648 69964 83700 69970
rect 83648 69906 83700 69912
rect 84200 69964 84252 69970
rect 84200 69906 84252 69912
rect 84936 69964 84988 69970
rect 84936 69906 84988 69912
rect 85488 69964 85540 69970
rect 85488 69906 85540 69912
rect 86132 69964 86184 69970
rect 86132 69906 86184 69912
rect 86776 69964 86828 69970
rect 86776 69906 86828 69912
rect 87420 69964 87472 69970
rect 87420 69906 87472 69912
rect 88064 69964 88116 69970
rect 88064 69906 88116 69912
rect 89352 69964 89404 69970
rect 89352 69906 89404 69912
rect 94688 69964 94740 69970
rect 94688 69906 94740 69912
rect 95792 69964 95844 69970
rect 95792 69906 95844 69912
rect 96436 69964 96488 69970
rect 96436 69906 96488 69912
rect 97080 69964 97132 69970
rect 97080 69906 97132 69912
rect 97724 69964 97776 69970
rect 97724 69906 97776 69912
rect 98368 69964 98420 69970
rect 98368 69906 98420 69912
rect 99012 69964 99064 69970
rect 99012 69906 99064 69912
rect 99656 69964 99708 69970
rect 99656 69906 99708 69912
rect 100300 69964 100352 69970
rect 100300 69906 100352 69912
rect 100944 69964 100996 69970
rect 100944 69906 100996 69912
rect 102140 69964 102192 69970
rect 102140 69906 102192 69912
rect 102232 69964 102284 69970
rect 102232 69906 102284 69912
rect 102876 69964 102928 69970
rect 102876 69906 102928 69912
rect 103152 69964 103204 69970
rect 103152 69906 103204 69912
rect 103520 69964 103572 69970
rect 103520 69906 103572 69912
rect 104624 69964 104676 69970
rect 104624 69906 104676 69912
rect 71976 68950 72004 69906
rect 71964 68944 72016 68950
rect 71964 68886 72016 68892
rect 72620 68406 72648 69906
rect 72608 68400 72660 68406
rect 72608 68342 72660 68348
rect 70492 68060 70544 68066
rect 70492 68002 70544 68008
rect 70398 67960 70454 67969
rect 70398 67895 70454 67904
rect 73356 65346 73384 69906
rect 73712 69896 73764 69902
rect 73712 69838 73764 69844
rect 73724 69562 73752 69838
rect 73712 69556 73764 69562
rect 73712 69498 73764 69504
rect 74000 66638 74028 69906
rect 74552 68241 74580 69906
rect 74538 68232 74594 68241
rect 74538 68167 74594 68176
rect 73988 66632 74040 66638
rect 73988 66574 74040 66580
rect 75196 65822 75224 69906
rect 75368 69828 75420 69834
rect 75368 69770 75420 69776
rect 75276 69760 75328 69766
rect 75276 69702 75328 69708
rect 75288 69630 75316 69702
rect 75380 69630 75408 69770
rect 75276 69624 75328 69630
rect 75276 69566 75328 69572
rect 75368 69624 75420 69630
rect 75368 69566 75420 69572
rect 76576 68678 76604 69906
rect 77128 68746 77156 69906
rect 77772 68882 77800 69906
rect 77760 68876 77812 68882
rect 77760 68818 77812 68824
rect 77772 68785 77800 68818
rect 77758 68776 77814 68785
rect 77116 68740 77168 68746
rect 77758 68711 77814 68720
rect 77116 68682 77168 68688
rect 76564 68672 76616 68678
rect 76564 68614 76616 68620
rect 78416 65929 78444 69906
rect 78402 65920 78458 65929
rect 78402 65855 78458 65864
rect 75184 65816 75236 65822
rect 75184 65758 75236 65764
rect 79060 65550 79088 69906
rect 79704 68377 79732 69906
rect 79690 68368 79746 68377
rect 79690 68303 79746 68312
rect 80440 67250 80468 69906
rect 81084 68542 81112 69906
rect 81072 68536 81124 68542
rect 81072 68478 81124 68484
rect 80428 67244 80480 67250
rect 80428 67186 80480 67192
rect 79048 65544 79100 65550
rect 79048 65486 79100 65492
rect 73344 65340 73396 65346
rect 73344 65282 73396 65288
rect 69848 64388 69900 64394
rect 69848 64330 69900 64336
rect 81728 64326 81756 69906
rect 82924 67182 82952 69906
rect 82912 67176 82964 67182
rect 82912 67118 82964 67124
rect 83660 66094 83688 69906
rect 84016 69828 84068 69834
rect 84016 69770 84068 69776
rect 84028 69630 84056 69770
rect 84016 69624 84068 69630
rect 84016 69566 84068 69572
rect 84212 68513 84240 69906
rect 84476 69896 84528 69902
rect 84476 69838 84528 69844
rect 84488 69562 84516 69838
rect 84476 69556 84528 69562
rect 84476 69498 84528 69504
rect 84198 68504 84254 68513
rect 84198 68439 84254 68448
rect 83648 66088 83700 66094
rect 83648 66030 83700 66036
rect 84948 65890 84976 69906
rect 85500 66230 85528 69906
rect 86144 68270 86172 69906
rect 86788 68474 86816 69906
rect 86776 68468 86828 68474
rect 86776 68410 86828 68416
rect 86132 68264 86184 68270
rect 86132 68206 86184 68212
rect 87432 68134 87460 69906
rect 87420 68128 87472 68134
rect 87420 68070 87472 68076
rect 88076 67153 88104 69906
rect 89364 68921 89392 69906
rect 89904 69896 89956 69902
rect 89904 69838 89956 69844
rect 89996 69896 90048 69902
rect 89996 69838 90048 69844
rect 90640 69896 90692 69902
rect 90640 69838 90692 69844
rect 91284 69896 91336 69902
rect 91284 69838 91336 69844
rect 91928 69896 91980 69902
rect 91928 69838 91980 69844
rect 92572 69896 92624 69902
rect 92572 69838 92624 69844
rect 93216 69896 93268 69902
rect 93216 69838 93268 69844
rect 93860 69896 93912 69902
rect 93860 69838 93912 69844
rect 89916 69630 89944 69838
rect 89904 69624 89956 69630
rect 89904 69566 89956 69572
rect 89350 68912 89406 68921
rect 89350 68847 89406 68856
rect 88062 67144 88118 67153
rect 88062 67079 88118 67088
rect 85488 66224 85540 66230
rect 85488 66166 85540 66172
rect 84936 65884 84988 65890
rect 84936 65826 84988 65832
rect 90008 65754 90036 69838
rect 89996 65748 90048 65754
rect 89996 65690 90048 65696
rect 90652 65278 90680 69838
rect 91296 66162 91324 69838
rect 91940 68882 91968 69838
rect 91928 68876 91980 68882
rect 91928 68818 91980 68824
rect 92584 68814 92612 69838
rect 92572 68808 92624 68814
rect 92572 68750 92624 68756
rect 93228 68610 93256 69838
rect 93216 68604 93268 68610
rect 93216 68546 93268 68552
rect 93872 67046 93900 69838
rect 93860 67040 93912 67046
rect 93860 66982 93912 66988
rect 91284 66156 91336 66162
rect 91284 66098 91336 66104
rect 94700 66026 94728 69906
rect 95148 68876 95200 68882
rect 95148 68818 95200 68824
rect 95160 68649 95188 68818
rect 95146 68640 95202 68649
rect 95146 68575 95202 68584
rect 95804 67114 95832 69906
rect 96448 68338 96476 69906
rect 97092 68882 97120 69906
rect 97736 69018 97764 69906
rect 97724 69012 97776 69018
rect 97724 68954 97776 68960
rect 97080 68876 97132 68882
rect 97080 68818 97132 68824
rect 96436 68332 96488 68338
rect 96436 68274 96488 68280
rect 95792 67108 95844 67114
rect 95792 67050 95844 67056
rect 98380 66842 98408 69906
rect 99024 66978 99052 69906
rect 99668 67522 99696 69906
rect 99656 67516 99708 67522
rect 99656 67458 99708 67464
rect 99012 66972 99064 66978
rect 99012 66914 99064 66920
rect 100312 66910 100340 69906
rect 100956 67425 100984 69906
rect 102152 69766 102180 69906
rect 102140 69760 102192 69766
rect 102140 69702 102192 69708
rect 100942 67416 100998 67425
rect 100942 67351 100998 67360
rect 100300 66904 100352 66910
rect 100300 66846 100352 66852
rect 98368 66836 98420 66842
rect 98368 66778 98420 66784
rect 94688 66020 94740 66026
rect 94688 65962 94740 65968
rect 102244 65618 102272 69906
rect 102888 67454 102916 69906
rect 103164 69630 103192 69906
rect 103152 69624 103204 69630
rect 103152 69566 103204 69572
rect 102876 67448 102928 67454
rect 102876 67390 102928 67396
rect 103532 66201 103560 69906
rect 104636 69154 104664 69906
rect 104624 69148 104676 69154
rect 104624 69090 104676 69096
rect 104164 69012 104216 69018
rect 104164 68954 104216 68960
rect 104176 68678 104204 68954
rect 104072 68672 104124 68678
rect 104072 68614 104124 68620
rect 104164 68672 104216 68678
rect 104164 68614 104216 68620
rect 104084 68490 104112 68614
rect 104084 68462 104296 68490
rect 104268 68338 104296 68462
rect 104164 68332 104216 68338
rect 104164 68274 104216 68280
rect 104256 68332 104308 68338
rect 104256 68274 104308 68280
rect 104176 67998 104204 68274
rect 104164 67992 104216 67998
rect 104164 67934 104216 67940
rect 106016 67590 106044 70722
rect 106004 67584 106056 67590
rect 106004 67526 106056 67532
rect 103980 67312 104032 67318
rect 104164 67312 104216 67318
rect 104032 67272 104164 67300
rect 103980 67254 104032 67260
rect 104164 67254 104216 67260
rect 106108 66706 106136 71538
rect 106200 70417 106228 71726
rect 106186 70408 106242 70417
rect 106186 70343 106242 70352
rect 106188 70304 106240 70310
rect 106188 70246 106240 70252
rect 106200 69086 106228 70246
rect 106188 69080 106240 69086
rect 106188 69022 106240 69028
rect 106292 68814 106320 198426
rect 107212 198422 107240 199786
rect 107488 198665 107516 199922
rect 108120 199708 108172 199714
rect 108120 199650 108172 199656
rect 107474 198656 107530 198665
rect 107474 198591 107530 198600
rect 106924 198416 106976 198422
rect 106924 198358 106976 198364
rect 107200 198416 107252 198422
rect 107200 198358 107252 198364
rect 106464 149116 106516 149122
rect 106464 149058 106516 149064
rect 106370 108488 106426 108497
rect 106370 108423 106426 108432
rect 106280 68808 106332 68814
rect 106280 68750 106332 68756
rect 106096 66700 106148 66706
rect 106096 66642 106148 66648
rect 103518 66192 103574 66201
rect 103518 66127 103574 66136
rect 106278 66056 106334 66065
rect 106278 65991 106334 66000
rect 102232 65612 102284 65618
rect 102232 65554 102284 65560
rect 106292 65346 106320 65991
rect 106280 65340 106332 65346
rect 106280 65282 106332 65288
rect 90640 65272 90692 65278
rect 90640 65214 90692 65220
rect 81716 64320 81768 64326
rect 81716 64262 81768 64268
rect 69388 64252 69440 64258
rect 69388 64194 69440 64200
rect 106384 20670 106412 108423
rect 106476 104825 106504 149058
rect 106462 104816 106518 104825
rect 106462 104751 106518 104760
rect 106462 102368 106518 102377
rect 106462 102303 106518 102312
rect 106476 69766 106504 102303
rect 106554 97880 106610 97889
rect 106554 97815 106610 97824
rect 106464 69760 106516 69766
rect 106464 69702 106516 69708
rect 106568 67318 106596 97815
rect 106936 78742 106964 198358
rect 107488 198150 107516 198591
rect 107476 198144 107528 198150
rect 107476 198086 107528 198092
rect 107014 169008 107070 169017
rect 107014 168943 107070 168952
rect 106924 78736 106976 78742
rect 106924 78678 106976 78684
rect 106556 67312 106608 67318
rect 106556 67254 106608 67260
rect 107028 66065 107056 168943
rect 107658 109032 107714 109041
rect 107658 108967 107660 108976
rect 107712 108967 107714 108976
rect 107660 108938 107712 108944
rect 108028 108928 108080 108934
rect 108028 108870 108080 108876
rect 108040 108497 108068 108870
rect 108026 108488 108082 108497
rect 108026 108423 108082 108432
rect 108028 104848 108080 104854
rect 108026 104816 108028 104825
rect 108080 104816 108082 104825
rect 108026 104751 108082 104760
rect 107660 99340 107712 99346
rect 107660 99282 107712 99288
rect 107672 98977 107700 99282
rect 107658 98968 107714 98977
rect 107658 98903 107714 98912
rect 107752 98660 107804 98666
rect 107752 98602 107804 98608
rect 107660 97980 107712 97986
rect 107660 97922 107712 97928
rect 107672 97617 107700 97922
rect 107764 97889 107792 98602
rect 107750 97880 107806 97889
rect 107750 97815 107806 97824
rect 107658 97608 107714 97617
rect 107658 97543 107714 97552
rect 107844 96620 107896 96626
rect 107844 96562 107896 96568
rect 107660 96552 107712 96558
rect 107660 96494 107712 96500
rect 107750 96520 107806 96529
rect 107672 96257 107700 96494
rect 107750 96455 107806 96464
rect 107658 96248 107714 96257
rect 107658 96183 107714 96192
rect 107764 95266 107792 96455
rect 107856 95577 107884 96562
rect 107842 95568 107898 95577
rect 107842 95503 107898 95512
rect 107752 95260 107804 95266
rect 107752 95202 107804 95208
rect 107660 95192 107712 95198
rect 107660 95134 107712 95140
rect 107672 94897 107700 95134
rect 107658 94888 107714 94897
rect 107658 94823 107714 94832
rect 107660 94512 107712 94518
rect 107660 94454 107712 94460
rect 107672 94217 107700 94454
rect 107658 94208 107714 94217
rect 107658 94143 107714 94152
rect 107752 93832 107804 93838
rect 107752 93774 107804 93780
rect 107660 93764 107712 93770
rect 107660 93706 107712 93712
rect 107672 93537 107700 93706
rect 107658 93528 107714 93537
rect 107658 93463 107714 93472
rect 107764 92857 107792 93774
rect 107750 92848 107806 92857
rect 107750 92783 107806 92792
rect 107752 91792 107804 91798
rect 107752 91734 107804 91740
rect 107764 91497 107792 91734
rect 107750 91488 107806 91497
rect 107750 91423 107806 91432
rect 107660 90364 107712 90370
rect 107660 90306 107712 90312
rect 107672 90137 107700 90306
rect 107658 90128 107714 90137
rect 107658 90063 107714 90072
rect 107108 89752 107160 89758
rect 107764 89714 107792 91423
rect 108026 90808 108082 90817
rect 108026 90743 108082 90752
rect 108040 90438 108068 90743
rect 108028 90432 108080 90438
rect 108028 90374 108080 90380
rect 107108 89694 107160 89700
rect 107120 69562 107148 89694
rect 107672 89686 107792 89714
rect 107292 88392 107344 88398
rect 107292 88334 107344 88340
rect 107200 85604 107252 85610
rect 107200 85546 107252 85552
rect 107108 69556 107160 69562
rect 107108 69498 107160 69504
rect 107014 66056 107070 66065
rect 107014 65991 107070 66000
rect 107212 65958 107240 85546
rect 107304 69834 107332 88334
rect 107384 81456 107436 81462
rect 107384 81398 107436 81404
rect 107292 69828 107344 69834
rect 107292 69770 107344 69776
rect 107396 66774 107424 81398
rect 107568 71800 107620 71806
rect 107568 71742 107620 71748
rect 107384 66768 107436 66774
rect 107384 66710 107436 66716
rect 107200 65952 107252 65958
rect 107200 65894 107252 65900
rect 107580 65793 107608 71742
rect 107566 65784 107622 65793
rect 107566 65719 107622 65728
rect 106372 20664 106424 20670
rect 106372 20606 106424 20612
rect 107672 4826 107700 89686
rect 107752 80028 107804 80034
rect 107752 79970 107804 79976
rect 107764 79937 107792 79970
rect 107750 79928 107806 79937
rect 107750 79863 107806 79872
rect 107936 78736 107988 78742
rect 107936 78678 107988 78684
rect 107752 78668 107804 78674
rect 107752 78610 107804 78616
rect 107764 77897 107792 78610
rect 107750 77888 107806 77897
rect 107750 77823 107806 77832
rect 107752 77240 107804 77246
rect 107750 77208 107752 77217
rect 107804 77208 107806 77217
rect 107750 77143 107806 77152
rect 107844 76016 107896 76022
rect 107750 75984 107806 75993
rect 107844 75958 107896 75964
rect 107750 75919 107752 75928
rect 107804 75919 107806 75928
rect 107752 75890 107804 75896
rect 107856 75857 107884 75958
rect 107842 75848 107898 75857
rect 107842 75783 107898 75792
rect 107844 75268 107896 75274
rect 107844 75210 107896 75216
rect 107752 75200 107804 75206
rect 107750 75168 107752 75177
rect 107804 75168 107806 75177
rect 107750 75103 107806 75112
rect 107752 74520 107804 74526
rect 107750 74488 107752 74497
rect 107804 74488 107806 74497
rect 107750 74423 107806 74432
rect 107752 73160 107804 73166
rect 107856 73137 107884 75210
rect 107752 73102 107804 73108
rect 107842 73128 107898 73137
rect 107764 72457 107792 73102
rect 107842 73063 107898 73072
rect 107750 72448 107806 72457
rect 107750 72383 107806 72392
rect 107948 65550 107976 78678
rect 108040 70378 108068 90374
rect 108132 76022 108160 199650
rect 108672 199640 108724 199646
rect 108672 199582 108724 199588
rect 108396 197872 108448 197878
rect 108396 197814 108448 197820
rect 108304 169584 108356 169590
rect 108304 169526 108356 169532
rect 108212 110560 108264 110566
rect 108212 110502 108264 110508
rect 108224 104417 108252 110502
rect 108210 104408 108266 104417
rect 108210 104343 108266 104352
rect 108212 103420 108264 103426
rect 108212 103362 108264 103368
rect 108224 102377 108252 103362
rect 108210 102368 108266 102377
rect 108210 102303 108266 102312
rect 108212 85536 108264 85542
rect 108212 85478 108264 85484
rect 108224 84697 108252 85478
rect 108210 84688 108266 84697
rect 108210 84623 108266 84632
rect 108316 84194 108344 169526
rect 108408 96694 108436 197814
rect 108578 196616 108634 196625
rect 108578 196551 108634 196560
rect 108488 193928 108540 193934
rect 108488 193870 108540 193876
rect 108500 165578 108528 193870
rect 108488 165572 108540 165578
rect 108488 165514 108540 165520
rect 108396 96688 108448 96694
rect 108396 96630 108448 96636
rect 108224 84166 108344 84194
rect 108120 76016 108172 76022
rect 108120 75958 108172 75964
rect 108224 75290 108252 84166
rect 108132 75262 108252 75290
rect 108028 70372 108080 70378
rect 108028 70314 108080 70320
rect 108132 68406 108160 75262
rect 108120 68400 108172 68406
rect 108120 68342 108172 68348
rect 108408 66230 108436 96630
rect 108500 87417 108528 165514
rect 108592 124370 108620 196551
rect 108580 124364 108632 124370
rect 108580 124306 108632 124312
rect 108592 110566 108620 124306
rect 108684 124302 108712 199582
rect 108776 198626 108804 199922
rect 108764 198620 108816 198626
rect 108764 198562 108816 198568
rect 109040 197940 109092 197946
rect 109040 197882 109092 197888
rect 108764 196784 108816 196790
rect 108764 196726 108816 196732
rect 108854 196752 108910 196761
rect 108776 165442 108804 196726
rect 108854 196687 108910 196696
rect 108868 165510 108896 196687
rect 108856 165504 108908 165510
rect 108856 165446 108908 165452
rect 108764 165436 108816 165442
rect 108764 165378 108816 165384
rect 108672 124296 108724 124302
rect 108672 124238 108724 124244
rect 108580 110560 108632 110566
rect 108580 110502 108632 110508
rect 108580 110356 108632 110362
rect 108580 110298 108632 110304
rect 108592 109857 108620 110298
rect 108578 109848 108634 109857
rect 108578 109783 108634 109792
rect 108580 101788 108632 101794
rect 108580 101730 108632 101736
rect 108592 89010 108620 101730
rect 108684 89457 108712 124238
rect 108776 101794 108804 165378
rect 108764 101788 108816 101794
rect 108764 101730 108816 101736
rect 108764 101652 108816 101658
rect 108764 101594 108816 101600
rect 108776 101017 108804 101594
rect 108762 101008 108818 101017
rect 108762 100943 108818 100952
rect 108764 100632 108816 100638
rect 108764 100574 108816 100580
rect 108776 99657 108804 100574
rect 108762 99648 108818 99657
rect 108762 99583 108818 99592
rect 108670 89448 108726 89457
rect 108670 89383 108726 89392
rect 108580 89004 108632 89010
rect 108580 88946 108632 88952
rect 108592 88777 108620 88946
rect 108578 88768 108634 88777
rect 108578 88703 108634 88712
rect 108486 87408 108542 87417
rect 108486 87343 108542 87352
rect 108500 71738 108528 87343
rect 108578 86048 108634 86057
rect 108578 85983 108634 85992
rect 108488 71732 108540 71738
rect 108488 71674 108540 71680
rect 108592 71670 108620 85983
rect 108868 82142 108896 165446
rect 108948 111784 109000 111790
rect 108948 111726 109000 111732
rect 108960 111217 108988 111726
rect 108946 111208 109002 111217
rect 108946 111143 109002 111152
rect 108948 110424 109000 110430
rect 108946 110392 108948 110401
rect 109000 110392 109002 110401
rect 108946 110327 109002 110336
rect 108948 107500 109000 107506
rect 108948 107442 109000 107448
rect 108960 107137 108988 107442
rect 108946 107128 109002 107137
rect 108946 107063 109002 107072
rect 108948 106684 109000 106690
rect 108948 106626 109000 106632
rect 108960 106457 108988 106626
rect 108946 106448 109002 106457
rect 108946 106383 109002 106392
rect 108948 106276 109000 106282
rect 108948 106218 109000 106224
rect 108960 105777 108988 106218
rect 108946 105768 109002 105777
rect 108946 105703 109002 105712
rect 108948 103488 109000 103494
rect 108948 103430 109000 103436
rect 108960 103057 108988 103430
rect 108946 103048 109002 103057
rect 108946 102983 109002 102992
rect 108948 102060 109000 102066
rect 108948 102002 109000 102008
rect 108960 101697 108988 102002
rect 108946 101688 109002 101697
rect 108946 101623 109002 101632
rect 108948 100700 109000 100706
rect 108948 100642 109000 100648
rect 108960 100337 108988 100642
rect 108946 100328 109002 100337
rect 108946 100263 109002 100272
rect 108948 88324 109000 88330
rect 108948 88266 109000 88272
rect 108960 88097 108988 88266
rect 108946 88088 109002 88097
rect 108946 88023 109002 88032
rect 108948 86964 109000 86970
rect 108948 86906 109000 86912
rect 108960 86737 108988 86906
rect 108946 86728 109002 86737
rect 108946 86663 109002 86672
rect 108948 84176 109000 84182
rect 108948 84118 109000 84124
rect 108960 84017 108988 84118
rect 108946 84008 109002 84017
rect 108946 83943 109002 83952
rect 108948 82816 109000 82822
rect 108948 82758 109000 82764
rect 108960 82657 108988 82758
rect 108946 82648 109002 82657
rect 108946 82583 109002 82592
rect 108856 82136 108908 82142
rect 108856 82078 108908 82084
rect 108868 81977 108896 82078
rect 108854 81968 108910 81977
rect 108854 81903 108910 81912
rect 108948 81388 109000 81394
rect 108948 81330 109000 81336
rect 108856 81320 108908 81326
rect 108854 81288 108856 81297
rect 108908 81288 108910 81297
rect 108854 81223 108910 81232
rect 108960 80617 108988 81330
rect 108946 80608 109002 80617
rect 108946 80543 109002 80552
rect 108672 79280 108724 79286
rect 108670 79248 108672 79257
rect 108724 79248 108726 79257
rect 108670 79183 108726 79192
rect 108580 71664 108632 71670
rect 108580 71606 108632 71612
rect 108684 70106 108712 79183
rect 108672 70100 108724 70106
rect 108672 70042 108724 70048
rect 109052 67318 109080 197882
rect 109132 197736 109184 197742
rect 109132 197678 109184 197684
rect 109144 68882 109172 197678
rect 109328 170542 109356 199922
rect 111156 199912 111208 199918
rect 111156 199854 111208 199860
rect 110420 198620 110472 198626
rect 110420 198562 110472 198568
rect 110236 188352 110288 188358
rect 110236 188294 110288 188300
rect 109316 170536 109368 170542
rect 109316 170478 109368 170484
rect 109224 170468 109276 170474
rect 109224 170410 109276 170416
rect 109236 169794 109264 170410
rect 109224 169788 109276 169794
rect 109224 169730 109276 169736
rect 109684 169788 109736 169794
rect 109684 169730 109736 169736
rect 109224 84856 109276 84862
rect 109224 84798 109276 84804
rect 109236 83337 109264 84798
rect 109222 83328 109278 83337
rect 109222 83263 109278 83272
rect 109132 68876 109184 68882
rect 109132 68818 109184 68824
rect 109040 67312 109092 67318
rect 109040 67254 109092 67260
rect 109696 67182 109724 169730
rect 110248 124166 110276 188294
rect 110328 183456 110380 183462
rect 110328 183398 110380 183404
rect 109776 124160 109828 124166
rect 109776 124102 109828 124108
rect 110236 124160 110288 124166
rect 110236 124102 110288 124108
rect 109788 122874 109816 124102
rect 109776 122868 109828 122874
rect 109776 122810 109828 122816
rect 109788 109002 109816 122810
rect 109776 108996 109828 109002
rect 109776 108938 109828 108944
rect 109774 87544 109830 87553
rect 109774 87479 109830 87488
rect 109040 67176 109092 67182
rect 109040 67118 109092 67124
rect 109684 67176 109736 67182
rect 109684 67118 109736 67124
rect 109052 66638 109080 67118
rect 109040 66632 109092 66638
rect 109040 66574 109092 66580
rect 108396 66224 108448 66230
rect 108396 66166 108448 66172
rect 107936 65544 107988 65550
rect 107936 65486 107988 65492
rect 109788 65414 109816 87479
rect 110340 70174 110368 183398
rect 110328 70168 110380 70174
rect 110328 70110 110380 70116
rect 110432 69034 110460 198562
rect 111064 198076 111116 198082
rect 111064 198018 111116 198024
rect 110512 197668 110564 197674
rect 110512 197610 110564 197616
rect 110340 69006 110460 69034
rect 110340 68762 110368 69006
rect 110340 68734 110460 68762
rect 110432 67522 110460 68734
rect 110524 67998 110552 197610
rect 110604 195492 110656 195498
rect 110604 195434 110656 195440
rect 110616 68610 110644 195434
rect 110696 169312 110748 169318
rect 110696 169254 110748 169260
rect 110708 168910 110736 169254
rect 110696 168904 110748 168910
rect 110696 168846 110748 168852
rect 111076 85678 111104 198018
rect 111168 197810 111196 199854
rect 111156 197804 111208 197810
rect 111156 197746 111208 197752
rect 111168 171902 111196 197746
rect 111260 174554 111288 199922
rect 112548 199782 112576 199922
rect 112536 199776 112588 199782
rect 112536 199718 112588 199724
rect 111800 198484 111852 198490
rect 111800 198426 111852 198432
rect 111248 174548 111300 174554
rect 111248 174490 111300 174496
rect 111156 171896 111208 171902
rect 111156 171838 111208 171844
rect 111156 168904 111208 168910
rect 111156 168846 111208 168852
rect 111064 85672 111116 85678
rect 111064 85614 111116 85620
rect 110604 68604 110656 68610
rect 110604 68546 110656 68552
rect 110512 67992 110564 67998
rect 110512 67934 110564 67940
rect 110420 67516 110472 67522
rect 110420 67458 110472 67464
rect 110524 67402 110552 67934
rect 110340 67374 110552 67402
rect 109776 65408 109828 65414
rect 109776 65350 109828 65356
rect 110340 64122 110368 67374
rect 110880 65816 110932 65822
rect 110880 65758 110932 65764
rect 110892 65414 110920 65758
rect 110880 65408 110932 65414
rect 110880 65350 110932 65356
rect 111076 64326 111104 85614
rect 111168 65822 111196 168846
rect 111248 167680 111300 167686
rect 111248 167622 111300 167628
rect 111260 68241 111288 167622
rect 111708 164960 111760 164966
rect 111708 164902 111760 164908
rect 111616 124908 111668 124914
rect 111616 124850 111668 124856
rect 111522 123448 111578 123457
rect 111522 123383 111578 123392
rect 111536 111790 111564 123383
rect 111524 111784 111576 111790
rect 111524 111726 111576 111732
rect 111628 77314 111656 124850
rect 111616 77308 111668 77314
rect 111616 77250 111668 77256
rect 111720 75206 111748 164902
rect 111708 75200 111760 75206
rect 111708 75142 111760 75148
rect 111812 68474 111840 198426
rect 111892 193860 111944 193866
rect 111892 193802 111944 193808
rect 111904 79286 111932 193802
rect 112444 181484 112496 181490
rect 112444 181426 112496 181432
rect 112456 180878 112484 181426
rect 112444 180872 112496 180878
rect 112444 180814 112496 180820
rect 111892 79280 111944 79286
rect 111892 79222 111944 79228
rect 111800 68468 111852 68474
rect 111800 68410 111852 68416
rect 112456 68338 112484 180814
rect 112548 171970 112576 199718
rect 113088 193996 113140 194002
rect 113088 193938 113140 193944
rect 112994 192536 113050 192545
rect 112994 192471 113050 192480
rect 112902 175944 112958 175953
rect 112902 175879 112958 175888
rect 112536 171964 112588 171970
rect 112536 171906 112588 171912
rect 112916 123486 112944 175879
rect 112536 123480 112588 123486
rect 112536 123422 112588 123428
rect 112904 123480 112956 123486
rect 112904 123422 112956 123428
rect 112548 81326 112576 123422
rect 113008 122942 113036 192471
rect 112996 122936 113048 122942
rect 112996 122878 113048 122884
rect 113008 106690 113036 122878
rect 112996 106684 113048 106690
rect 112996 106626 113048 106632
rect 112536 81320 112588 81326
rect 112536 81262 112588 81268
rect 113100 73817 113128 193938
rect 113086 73808 113142 73817
rect 113086 73743 113142 73752
rect 113086 71088 113142 71097
rect 113086 71023 113142 71032
rect 112444 68332 112496 68338
rect 112444 68274 112496 68280
rect 111246 68232 111302 68241
rect 111246 68167 111302 68176
rect 113100 67590 113128 71023
rect 113192 69154 113220 199922
rect 113824 199776 113876 199782
rect 113824 199718 113876 199724
rect 113732 199368 113784 199374
rect 113732 199310 113784 199316
rect 113744 198642 113772 199310
rect 113836 199306 113864 199718
rect 113824 199300 113876 199306
rect 113824 199242 113876 199248
rect 113744 198614 113864 198642
rect 113836 198558 113864 198614
rect 113824 198552 113876 198558
rect 113824 198494 113876 198500
rect 113272 195560 113324 195566
rect 113272 195502 113324 195508
rect 113180 69148 113232 69154
rect 113180 69090 113232 69096
rect 113284 68678 113312 195502
rect 113364 195424 113416 195430
rect 113364 195366 113416 195372
rect 113272 68672 113324 68678
rect 113376 68649 113404 195366
rect 113836 190534 113864 198494
rect 114480 198082 114508 199922
rect 114468 198076 114520 198082
rect 114468 198018 114520 198024
rect 114560 195288 114612 195294
rect 114560 195230 114612 195236
rect 113824 190528 113876 190534
rect 113824 190470 113876 190476
rect 113546 69456 113602 69465
rect 113546 69391 113602 69400
rect 113560 69154 113588 69391
rect 113836 69329 113864 190470
rect 114468 173256 114520 173262
rect 114468 173198 114520 173204
rect 114480 172582 114508 173198
rect 113916 172576 113968 172582
rect 113916 172518 113968 172524
rect 114468 172576 114520 172582
rect 114468 172518 114520 172524
rect 113822 69320 113878 69329
rect 113822 69255 113878 69264
rect 113548 69148 113600 69154
rect 113548 69090 113600 69096
rect 113272 68614 113324 68620
rect 113362 68640 113418 68649
rect 113362 68575 113418 68584
rect 113088 67584 113140 67590
rect 113088 67526 113140 67532
rect 113928 65929 113956 172518
rect 114572 93854 114600 195230
rect 115308 183462 115336 199922
rect 115664 194948 115716 194954
rect 115664 194890 115716 194896
rect 115296 183456 115348 183462
rect 115296 183398 115348 183404
rect 115308 169658 115336 183398
rect 115388 170604 115440 170610
rect 115388 170546 115440 170552
rect 115400 169862 115428 170546
rect 115388 169856 115440 169862
rect 115388 169798 115440 169804
rect 115296 169652 115348 169658
rect 115296 169594 115348 169600
rect 115400 161474 115428 169798
rect 115216 161446 115428 161474
rect 114572 93826 114692 93854
rect 114664 68513 114692 93826
rect 114650 68504 114706 68513
rect 114650 68439 114706 68448
rect 115216 67386 115244 161446
rect 115676 132494 115704 194890
rect 115756 193724 115808 193730
rect 115756 193666 115808 193672
rect 115308 132466 115704 132494
rect 115308 124438 115336 132466
rect 115296 124432 115348 124438
rect 115296 124374 115348 124380
rect 115308 102066 115336 124374
rect 115768 123010 115796 193666
rect 115860 190602 115888 199922
rect 115940 195356 115992 195362
rect 115940 195298 115992 195304
rect 115848 190596 115900 190602
rect 115848 190538 115900 190544
rect 115756 123004 115808 123010
rect 115756 122946 115808 122952
rect 115768 122834 115796 122946
rect 115400 122806 115796 122834
rect 115296 102060 115348 102066
rect 115296 102002 115348 102008
rect 115400 101658 115428 122806
rect 115388 101652 115440 101658
rect 115388 101594 115440 101600
rect 115860 74534 115888 190538
rect 115768 74506 115888 74534
rect 115768 70038 115796 74506
rect 115756 70032 115808 70038
rect 115756 69974 115808 69980
rect 115768 69086 115796 69974
rect 115756 69080 115808 69086
rect 115756 69022 115808 69028
rect 115952 68921 115980 195298
rect 116596 194682 116624 199922
rect 117136 198960 117188 198966
rect 117136 198902 117188 198908
rect 117044 198824 117096 198830
rect 117044 198766 117096 198772
rect 116584 194676 116636 194682
rect 116584 194618 116636 194624
rect 116596 71097 116624 194618
rect 116676 184204 116728 184210
rect 116676 184146 116728 184152
rect 116688 183598 116716 184146
rect 116676 183592 116728 183598
rect 116676 183534 116728 183540
rect 116582 71088 116638 71097
rect 116582 71023 116638 71032
rect 115938 68912 115994 68921
rect 115938 68847 115994 68856
rect 115846 68504 115902 68513
rect 115846 68439 115902 68448
rect 115860 68105 115888 68439
rect 116688 68377 116716 183534
rect 117056 124545 117084 198766
rect 117042 124536 117098 124545
rect 117042 124471 117098 124480
rect 117056 122834 117084 124471
rect 116872 122806 117084 122834
rect 116768 121508 116820 121514
rect 116768 121450 116820 121456
rect 116780 81394 116808 121450
rect 116872 109002 116900 122806
rect 117148 122126 117176 198902
rect 117228 198892 117280 198898
rect 117228 198834 117280 198840
rect 117136 122120 117188 122126
rect 117136 122062 117188 122068
rect 117148 121514 117176 122062
rect 117136 121508 117188 121514
rect 117136 121450 117188 121456
rect 116860 108996 116912 109002
rect 116860 108938 116912 108944
rect 117240 82890 117268 198834
rect 117332 198558 117360 199922
rect 117700 199238 117728 199922
rect 117688 199232 117740 199238
rect 117688 199174 117740 199180
rect 118516 198756 118568 198762
rect 118516 198698 118568 198704
rect 117320 198552 117372 198558
rect 117320 198494 117372 198500
rect 117964 197464 118016 197470
rect 117964 197406 118016 197412
rect 117976 194614 118004 197406
rect 117964 194608 118016 194614
rect 117964 194550 118016 194556
rect 117976 183462 118004 194550
rect 118056 190528 118108 190534
rect 118056 190470 118108 190476
rect 117964 183456 118016 183462
rect 117964 183398 118016 183404
rect 117228 82884 117280 82890
rect 117228 82826 117280 82832
rect 116768 81388 116820 81394
rect 116768 81330 116820 81336
rect 117976 73370 118004 183398
rect 118068 169454 118096 190470
rect 118056 169448 118108 169454
rect 118056 169390 118108 169396
rect 118528 78810 118556 198698
rect 118608 197396 118660 197402
rect 118608 197338 118660 197344
rect 118148 78804 118200 78810
rect 118148 78746 118200 78752
rect 118516 78804 118568 78810
rect 118516 78746 118568 78752
rect 118160 78674 118188 78746
rect 118148 78668 118200 78674
rect 118148 78610 118200 78616
rect 118620 76090 118648 197338
rect 118700 196036 118752 196042
rect 118700 195978 118752 195984
rect 118712 194002 118740 195978
rect 118700 193996 118752 194002
rect 118700 193938 118752 193944
rect 119080 130286 119108 200058
rect 119172 197470 119200 200246
rect 119160 197464 119212 197470
rect 119160 197406 119212 197412
rect 119264 195974 119292 209746
rect 119448 196790 119476 209746
rect 119804 204332 119856 204338
rect 119804 204274 119856 204280
rect 119632 197402 119660 200260
rect 119710 199472 119766 199481
rect 119710 199407 119766 199416
rect 119620 197396 119672 197402
rect 119620 197338 119672 197344
rect 119436 196784 119488 196790
rect 119436 196726 119488 196732
rect 119724 196042 119752 199407
rect 119712 196036 119764 196042
rect 119712 195978 119764 195984
rect 119172 195946 119292 195974
rect 119068 130280 119120 130286
rect 119068 130222 119120 130228
rect 119172 124166 119200 195946
rect 119342 165608 119398 165617
rect 119342 165543 119398 165552
rect 119356 164898 119384 165543
rect 119344 164892 119396 164898
rect 119344 164834 119396 164840
rect 119250 125488 119306 125497
rect 119250 125423 119306 125432
rect 119264 124642 119292 125423
rect 119252 124636 119304 124642
rect 119252 124578 119304 124584
rect 119160 124160 119212 124166
rect 119160 124102 119212 124108
rect 119264 96558 119292 124578
rect 119252 96552 119304 96558
rect 119252 96494 119304 96500
rect 119356 90370 119384 164834
rect 119816 132494 119844 204274
rect 119448 132466 119844 132494
rect 119448 123146 119476 132466
rect 119620 130280 119672 130286
rect 119620 130222 119672 130228
rect 119528 124160 119580 124166
rect 119528 124102 119580 124108
rect 119540 123282 119568 124102
rect 119528 123276 119580 123282
rect 119528 123218 119580 123224
rect 119436 123140 119488 123146
rect 119436 123082 119488 123088
rect 119344 90364 119396 90370
rect 119344 90306 119396 90312
rect 119448 86970 119476 123082
rect 119540 88330 119568 123218
rect 119632 98666 119660 130222
rect 119710 125352 119766 125361
rect 119710 125287 119766 125296
rect 119724 124506 119752 125287
rect 119908 124846 119936 224946
rect 120184 219881 120212 260102
rect 120356 258732 120408 258738
rect 120356 258674 120408 258680
rect 120170 219872 120226 219881
rect 120170 219807 120226 219816
rect 120170 217696 120226 217705
rect 120170 217631 120226 217640
rect 119988 212900 120040 212906
rect 119988 212842 120040 212848
rect 119896 124840 119948 124846
rect 119896 124782 119948 124788
rect 119712 124500 119764 124506
rect 119712 124442 119764 124448
rect 119620 98660 119672 98666
rect 119620 98602 119672 98608
rect 119724 96626 119752 124442
rect 119908 104854 119936 124782
rect 120000 111722 120028 212842
rect 120078 203416 120134 203425
rect 120078 203351 120134 203360
rect 120092 199714 120120 203351
rect 120080 199708 120132 199714
rect 120080 199650 120132 199656
rect 120184 193934 120212 217631
rect 120368 201385 120396 258674
rect 120448 220788 120500 220794
rect 120448 220730 120500 220736
rect 120460 220425 120488 220730
rect 120446 220416 120502 220425
rect 120446 220351 120502 220360
rect 120354 201376 120410 201385
rect 120354 201311 120410 201320
rect 120460 199646 120488 220351
rect 120736 218142 120764 700266
rect 121460 553444 121512 553450
rect 121460 553386 121512 553392
rect 120816 527196 120868 527202
rect 120816 527138 120868 527144
rect 120724 218136 120776 218142
rect 120724 218078 120776 218084
rect 120828 214062 120856 527138
rect 120908 253156 120960 253162
rect 120908 253098 120960 253104
rect 120920 229838 120948 253098
rect 121000 252680 121052 252686
rect 121000 252622 121052 252628
rect 121012 232694 121040 252622
rect 121368 252068 121420 252074
rect 121368 252010 121420 252016
rect 121276 251388 121328 251394
rect 121276 251330 121328 251336
rect 121092 250436 121144 250442
rect 121092 250378 121144 250384
rect 121104 233170 121132 250378
rect 121184 250028 121236 250034
rect 121184 249970 121236 249976
rect 121092 233164 121144 233170
rect 121092 233106 121144 233112
rect 121196 232830 121224 249970
rect 121288 245002 121316 251330
rect 121380 246498 121408 252010
rect 121472 248402 121500 553386
rect 121920 257372 121972 257378
rect 121920 257314 121972 257320
rect 121736 256012 121788 256018
rect 121736 255954 121788 255960
rect 121552 249144 121604 249150
rect 121552 249086 121604 249092
rect 121460 248396 121512 248402
rect 121460 248338 121512 248344
rect 121458 248296 121514 248305
rect 121458 248231 121514 248240
rect 121472 247110 121500 248231
rect 121460 247104 121512 247110
rect 121460 247046 121512 247052
rect 121458 246936 121514 246945
rect 121458 246871 121514 246880
rect 121368 246492 121420 246498
rect 121368 246434 121420 246440
rect 121472 245682 121500 246871
rect 121460 245676 121512 245682
rect 121460 245618 121512 245624
rect 121276 244996 121328 245002
rect 121276 244938 121328 244944
rect 121460 244452 121512 244458
rect 121460 244394 121512 244400
rect 121472 244361 121500 244394
rect 121458 244352 121514 244361
rect 121458 244287 121514 244296
rect 121564 242962 121592 249086
rect 121642 244896 121698 244905
rect 121642 244831 121698 244840
rect 121656 244390 121684 244831
rect 121644 244384 121696 244390
rect 121644 244326 121696 244332
rect 121552 242956 121604 242962
rect 121552 242898 121604 242904
rect 121458 242176 121514 242185
rect 121458 242111 121514 242120
rect 121472 241534 121500 242111
rect 121550 241632 121606 241641
rect 121550 241567 121552 241576
rect 121604 241567 121606 241576
rect 121552 241538 121604 241544
rect 121460 241528 121512 241534
rect 121460 241470 121512 241476
rect 121458 238096 121514 238105
rect 121458 238031 121514 238040
rect 121472 237402 121500 238031
rect 121380 237386 121500 237402
rect 121368 237380 121500 237386
rect 121420 237374 121500 237380
rect 121368 237322 121420 237328
rect 121276 233232 121328 233238
rect 121276 233174 121328 233180
rect 121184 232824 121236 232830
rect 121184 232766 121236 232772
rect 121000 232688 121052 232694
rect 121000 232630 121052 232636
rect 120908 229832 120960 229838
rect 120908 229774 120960 229780
rect 121000 218068 121052 218074
rect 121000 218010 121052 218016
rect 120816 214056 120868 214062
rect 120816 213998 120868 214004
rect 120722 208176 120778 208185
rect 120722 208111 120778 208120
rect 120448 199640 120500 199646
rect 120448 199582 120500 199588
rect 120172 193928 120224 193934
rect 120172 193870 120224 193876
rect 120630 166968 120686 166977
rect 120630 166903 120686 166912
rect 119988 111716 120040 111722
rect 119988 111658 120040 111664
rect 119896 104848 119948 104854
rect 119896 104790 119948 104796
rect 119712 96620 119764 96626
rect 119712 96562 119764 96568
rect 119986 95296 120042 95305
rect 119986 95231 120042 95240
rect 120000 94518 120028 95231
rect 120644 95198 120672 166903
rect 120736 120902 120764 208111
rect 121012 165374 121040 218010
rect 121184 212492 121236 212498
rect 121184 212434 121236 212440
rect 121092 205692 121144 205698
rect 121092 205634 121144 205640
rect 121000 165368 121052 165374
rect 121000 165310 121052 165316
rect 121012 161474 121040 165310
rect 120828 161446 121040 161474
rect 120724 120896 120776 120902
rect 120724 120838 120776 120844
rect 120080 95192 120132 95198
rect 120080 95134 120132 95140
rect 120632 95192 120684 95198
rect 120632 95134 120684 95140
rect 120092 94586 120120 95134
rect 120080 94580 120132 94586
rect 120080 94522 120132 94528
rect 119988 94512 120040 94518
rect 119988 94454 120040 94460
rect 119528 88324 119580 88330
rect 119528 88266 119580 88272
rect 119436 86964 119488 86970
rect 119436 86906 119488 86912
rect 120736 80034 120764 120838
rect 120828 90438 120856 161446
rect 121104 124710 121132 205634
rect 121092 124704 121144 124710
rect 121092 124646 121144 124652
rect 120908 124160 120960 124166
rect 120908 124102 120960 124108
rect 120920 123214 120948 124102
rect 120908 123208 120960 123214
rect 120908 123150 120960 123156
rect 120920 93770 120948 123150
rect 121104 97986 121132 124646
rect 121196 124166 121224 212434
rect 121288 124574 121316 233174
rect 121380 124778 121408 237322
rect 121460 230852 121512 230858
rect 121460 230794 121512 230800
rect 121472 230761 121500 230794
rect 121458 230752 121514 230761
rect 121458 230687 121514 230696
rect 121458 229256 121514 229265
rect 121458 229191 121514 229200
rect 121472 229158 121500 229191
rect 121460 229152 121512 229158
rect 121460 229094 121512 229100
rect 121564 225010 121592 241538
rect 121552 225004 121604 225010
rect 121552 224946 121604 224952
rect 121460 224936 121512 224942
rect 121460 224878 121512 224884
rect 121472 224641 121500 224878
rect 121458 224632 121514 224641
rect 121458 224567 121514 224576
rect 121550 222592 121606 222601
rect 121550 222527 121606 222536
rect 121460 222080 121512 222086
rect 121460 222022 121512 222028
rect 121472 221921 121500 222022
rect 121458 221912 121514 221921
rect 121458 221847 121514 221856
rect 121564 219434 121592 222527
rect 121472 219406 121592 219434
rect 121472 218074 121500 219406
rect 121552 218136 121604 218142
rect 121552 218078 121604 218084
rect 121460 218068 121512 218074
rect 121460 218010 121512 218016
rect 121564 217954 121592 218078
rect 121472 217926 121592 217954
rect 121472 216034 121500 217926
rect 121460 216028 121512 216034
rect 121460 215970 121512 215976
rect 121472 215801 121500 215970
rect 121458 215792 121514 215801
rect 121458 215727 121514 215736
rect 121458 214976 121514 214985
rect 121458 214911 121514 214920
rect 121472 213994 121500 214911
rect 121552 214056 121604 214062
rect 121552 213998 121604 214004
rect 121460 213988 121512 213994
rect 121460 213930 121512 213936
rect 121458 212256 121514 212265
rect 121458 212191 121514 212200
rect 121472 211818 121500 212191
rect 121460 211812 121512 211818
rect 121460 211754 121512 211760
rect 121460 211676 121512 211682
rect 121460 211618 121512 211624
rect 121472 204338 121500 211618
rect 121564 211041 121592 213998
rect 121550 211032 121606 211041
rect 121550 210967 121606 210976
rect 121550 206816 121606 206825
rect 121550 206751 121606 206760
rect 121564 206378 121592 206751
rect 121552 206372 121604 206378
rect 121552 206314 121604 206320
rect 121550 206136 121606 206145
rect 121550 206071 121606 206080
rect 121460 204332 121512 204338
rect 121460 204274 121512 204280
rect 121564 198762 121592 206071
rect 121656 198830 121684 244326
rect 121748 232801 121776 255954
rect 121828 248396 121880 248402
rect 121828 248338 121880 248344
rect 121840 239601 121868 248338
rect 121826 239592 121882 239601
rect 121826 239527 121882 239536
rect 121840 239494 121868 239527
rect 121828 239488 121880 239494
rect 121828 239430 121880 239436
rect 121828 237516 121880 237522
rect 121828 237458 121880 237464
rect 121840 237425 121868 237458
rect 121826 237416 121882 237425
rect 121826 237351 121882 237360
rect 121734 232792 121790 232801
rect 121734 232727 121790 232736
rect 121748 230926 121776 232727
rect 121736 230920 121788 230926
rect 121736 230862 121788 230868
rect 121736 213920 121788 213926
rect 121736 213862 121788 213868
rect 121748 213081 121776 213862
rect 121734 213072 121790 213081
rect 121734 213007 121790 213016
rect 121840 209774 121868 237351
rect 121932 222601 121960 257314
rect 122104 251932 122156 251938
rect 122104 251874 122156 251880
rect 122012 246356 122064 246362
rect 122012 246298 122064 246304
rect 122024 246265 122052 246298
rect 122010 246256 122066 246265
rect 122010 246191 122066 246200
rect 122012 245676 122064 245682
rect 122012 245618 122064 245624
rect 122024 233238 122052 245618
rect 122116 244934 122144 251874
rect 122196 251524 122248 251530
rect 122196 251466 122248 251472
rect 122208 246430 122236 251466
rect 122378 248976 122434 248985
rect 122378 248911 122434 248920
rect 122196 246424 122248 246430
rect 122196 246366 122248 246372
rect 122392 246362 122420 248911
rect 122380 246356 122432 246362
rect 122380 246298 122432 246304
rect 122654 245848 122710 245857
rect 122654 245783 122710 245792
rect 122668 245750 122696 245783
rect 122656 245744 122708 245750
rect 122656 245686 122708 245692
rect 122104 244928 122156 244934
rect 122104 244870 122156 244876
rect 122288 243024 122340 243030
rect 122286 242992 122288 243001
rect 122340 242992 122342 243001
rect 122104 242956 122156 242962
rect 122286 242927 122342 242936
rect 122104 242898 122156 242904
rect 122012 233232 122064 233238
rect 122012 233174 122064 233180
rect 121918 222592 121974 222601
rect 121918 222527 121974 222536
rect 122012 217320 122064 217326
rect 122012 217262 122064 217268
rect 122024 217025 122052 217262
rect 122010 217016 122066 217025
rect 122010 216951 122066 216960
rect 121918 213616 121974 213625
rect 121918 213551 121974 213560
rect 121932 212566 121960 213551
rect 121920 212560 121972 212566
rect 121920 212502 121972 212508
rect 122024 212378 122052 216951
rect 122116 212906 122144 242898
rect 122286 235376 122342 235385
rect 122286 235311 122342 235320
rect 122300 234734 122328 235311
rect 122288 234728 122340 234734
rect 122288 234670 122340 234676
rect 122470 234696 122526 234705
rect 122470 234631 122472 234640
rect 122524 234631 122526 234640
rect 122472 234602 122524 234608
rect 122470 233336 122526 233345
rect 122470 233271 122472 233280
rect 122524 233271 122526 233280
rect 122472 233242 122524 233248
rect 122288 230920 122340 230926
rect 122288 230862 122340 230868
rect 122194 223816 122250 223825
rect 122194 223751 122250 223760
rect 122104 212900 122156 212906
rect 122104 212842 122156 212848
rect 121932 212350 122052 212378
rect 121932 211682 121960 212350
rect 122012 211812 122064 211818
rect 122012 211754 122064 211760
rect 121920 211676 121972 211682
rect 121920 211618 121972 211624
rect 121840 209746 121960 209774
rect 121734 205456 121790 205465
rect 121734 205391 121790 205400
rect 121644 198824 121696 198830
rect 121644 198766 121696 198772
rect 121552 198756 121604 198762
rect 121552 198698 121604 198704
rect 121748 195974 121776 205391
rect 121826 202056 121882 202065
rect 121826 201991 121882 202000
rect 121840 201550 121868 201991
rect 121828 201544 121880 201550
rect 121828 201486 121880 201492
rect 121472 195946 121776 195974
rect 121472 124914 121500 195946
rect 121932 194954 121960 209746
rect 122024 198898 122052 211754
rect 122104 206372 122156 206378
rect 122104 206314 122156 206320
rect 122012 198892 122064 198898
rect 122012 198834 122064 198840
rect 121920 194948 121972 194954
rect 121920 194890 121972 194896
rect 122116 193866 122144 206314
rect 122104 193860 122156 193866
rect 122104 193802 122156 193808
rect 122104 169176 122156 169182
rect 122104 169118 122156 169124
rect 121460 124908 121512 124914
rect 121460 124850 121512 124856
rect 121368 124772 121420 124778
rect 121368 124714 121420 124720
rect 121276 124568 121328 124574
rect 121276 124510 121328 124516
rect 121184 124160 121236 124166
rect 121184 124102 121236 124108
rect 121288 110362 121316 124510
rect 121276 110356 121328 110362
rect 121276 110298 121328 110304
rect 121380 103426 121408 124714
rect 121368 103420 121420 103426
rect 121368 103362 121420 103368
rect 121092 97980 121144 97986
rect 121092 97922 121144 97928
rect 120908 93764 120960 93770
rect 120908 93706 120960 93712
rect 120816 90432 120868 90438
rect 120816 90374 120868 90380
rect 120724 80028 120776 80034
rect 120724 79970 120776 79976
rect 118148 76084 118200 76090
rect 118148 76026 118200 76032
rect 118608 76084 118660 76090
rect 118608 76026 118660 76032
rect 118160 75274 118188 76026
rect 118148 75268 118200 75274
rect 118148 75210 118200 75216
rect 117964 73364 118016 73370
rect 117964 73306 118016 73312
rect 117976 73166 118004 73306
rect 117964 73160 118016 73166
rect 117964 73102 118016 73108
rect 117226 68912 117282 68921
rect 117226 68847 117282 68856
rect 117240 68513 117268 68847
rect 117226 68504 117282 68513
rect 117226 68439 117282 68448
rect 116674 68368 116730 68377
rect 116674 68303 116730 68312
rect 115846 68096 115902 68105
rect 115846 68031 115902 68040
rect 115204 67380 115256 67386
rect 115204 67322 115256 67328
rect 115848 67380 115900 67386
rect 115848 67322 115900 67328
rect 115860 66774 115888 67322
rect 115848 66768 115900 66774
rect 115848 66710 115900 66716
rect 121460 66088 121512 66094
rect 121460 66030 121512 66036
rect 113914 65920 113970 65929
rect 113914 65855 113970 65864
rect 121472 65822 121500 66030
rect 122116 65822 122144 169118
rect 122208 132494 122236 223751
rect 122300 205698 122328 230862
rect 122470 225856 122526 225865
rect 122470 225791 122526 225800
rect 122484 225622 122512 225791
rect 122472 225616 122524 225622
rect 122472 225558 122524 225564
rect 122484 212498 122512 225558
rect 122472 212492 122524 212498
rect 122472 212434 122524 212440
rect 122378 208856 122434 208865
rect 122378 208791 122434 208800
rect 122288 205692 122340 205698
rect 122288 205634 122340 205640
rect 122392 198966 122420 208791
rect 122562 205456 122618 205465
rect 122562 205391 122618 205400
rect 122576 204950 122604 205391
rect 122564 204944 122616 204950
rect 122564 204886 122616 204892
rect 122562 204096 122618 204105
rect 122562 204031 122618 204040
rect 122576 202910 122604 204031
rect 122564 202904 122616 202910
rect 122564 202846 122616 202852
rect 122562 201376 122618 201385
rect 122562 201311 122618 201320
rect 122576 200190 122604 201311
rect 122564 200184 122616 200190
rect 122564 200126 122616 200132
rect 122380 198960 122432 198966
rect 122380 198902 122432 198908
rect 122668 188358 122696 245686
rect 122746 236056 122802 236065
rect 122746 235991 122748 236000
rect 122800 235991 122802 236000
rect 122748 235962 122800 235968
rect 122760 193730 122788 235962
rect 122852 198529 122880 700402
rect 137848 700398 137876 703520
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 153212 702406 154160 702434
rect 169772 702406 170352 702434
rect 137836 700392 137888 700398
rect 137836 700334 137888 700340
rect 123668 265668 123720 265674
rect 123668 265610 123720 265616
rect 123574 252784 123630 252793
rect 123574 252719 123630 252728
rect 123484 249960 123536 249966
rect 123484 249902 123536 249908
rect 123496 206310 123524 249902
rect 123588 209778 123616 252719
rect 123680 222086 123708 265610
rect 126336 254584 126388 254590
rect 126336 254526 126388 254532
rect 142896 254584 142948 254590
rect 142896 254526 142948 254532
rect 124864 253496 124916 253502
rect 124864 253438 124916 253444
rect 124036 253020 124088 253026
rect 124036 252962 124088 252968
rect 123758 252648 123814 252657
rect 123758 252583 123814 252592
rect 123668 222080 123720 222086
rect 123668 222022 123720 222028
rect 123772 215966 123800 252583
rect 123852 250708 123904 250714
rect 123852 250650 123904 250656
rect 123760 215960 123812 215966
rect 123760 215902 123812 215908
rect 123864 214606 123892 250650
rect 123944 250368 123996 250374
rect 123944 250310 123996 250316
rect 123956 214674 123984 250310
rect 124048 224874 124076 252962
rect 124220 252136 124272 252142
rect 124220 252078 124272 252084
rect 124128 251592 124180 251598
rect 124128 251534 124180 251540
rect 124140 239426 124168 251534
rect 124128 239420 124180 239426
rect 124128 239362 124180 239368
rect 124036 224868 124088 224874
rect 124036 224810 124088 224816
rect 123944 214668 123996 214674
rect 123944 214610 123996 214616
rect 123852 214600 123904 214606
rect 123852 214542 123904 214548
rect 123576 209772 123628 209778
rect 123576 209714 123628 209720
rect 123484 206304 123536 206310
rect 123484 206246 123536 206252
rect 122838 198520 122894 198529
rect 122838 198455 122894 198464
rect 122748 193724 122800 193730
rect 122748 193666 122800 193672
rect 123484 189848 123536 189854
rect 123484 189790 123536 189796
rect 123496 189106 123524 189790
rect 123484 189100 123536 189106
rect 123484 189042 123536 189048
rect 122656 188352 122708 188358
rect 122656 188294 122708 188300
rect 123496 183002 123524 189042
rect 123852 183456 123904 183462
rect 123852 183398 123904 183404
rect 123404 182974 123524 183002
rect 123404 180794 123432 182974
rect 123484 182844 123536 182850
rect 123484 182786 123536 182792
rect 123496 182238 123524 182786
rect 123484 182232 123536 182238
rect 123484 182174 123536 182180
rect 123496 181914 123524 182174
rect 123496 181886 123616 181914
rect 123404 180766 123524 180794
rect 123208 177404 123260 177410
rect 123208 177346 123260 177352
rect 123220 176730 123248 177346
rect 123208 176724 123260 176730
rect 123208 176666 123260 176672
rect 122208 132466 122328 132494
rect 122300 129062 122328 132466
rect 122288 129056 122340 129062
rect 122288 128998 122340 129004
rect 122194 122904 122250 122913
rect 122194 122839 122250 122848
rect 122208 84862 122236 122839
rect 122300 91798 122328 128998
rect 122288 91792 122340 91798
rect 122288 91734 122340 91740
rect 122196 84856 122248 84862
rect 122196 84798 122248 84804
rect 123496 65890 123524 180766
rect 123588 68270 123616 181886
rect 123668 176724 123720 176730
rect 123668 176666 123720 176672
rect 123576 68264 123628 68270
rect 123576 68206 123628 68212
rect 123680 66162 123708 176666
rect 123760 171964 123812 171970
rect 123760 171906 123812 171912
rect 123772 171154 123800 171906
rect 123760 171148 123812 171154
rect 123760 171090 123812 171096
rect 123772 67386 123800 171090
rect 123864 168298 123892 183398
rect 123852 168292 123904 168298
rect 123852 168234 123904 168240
rect 124232 114442 124260 252078
rect 124312 251796 124364 251802
rect 124312 251738 124364 251744
rect 124324 114510 124352 251738
rect 124876 207670 124904 253438
rect 126244 253292 126296 253298
rect 126244 253234 126296 253240
rect 125140 251728 125192 251734
rect 125140 251670 125192 251676
rect 125048 250776 125100 250782
rect 125048 250718 125100 250724
rect 124956 250300 125008 250306
rect 124956 250242 125008 250248
rect 124968 221474 124996 250242
rect 125060 229090 125088 250718
rect 125152 240786 125180 251670
rect 125140 240780 125192 240786
rect 125140 240722 125192 240728
rect 125048 229084 125100 229090
rect 125048 229026 125100 229032
rect 125048 222216 125100 222222
rect 125048 222158 125100 222164
rect 124956 221468 125008 221474
rect 124956 221410 125008 221416
rect 124864 207664 124916 207670
rect 124864 207606 124916 207612
rect 124404 201544 124456 201550
rect 124404 201486 124456 201492
rect 124416 165306 124444 201486
rect 125060 199782 125088 222158
rect 125048 199776 125100 199782
rect 125048 199718 125100 199724
rect 125600 170672 125652 170678
rect 125600 170614 125652 170620
rect 124404 165300 124456 165306
rect 124404 165242 124456 165248
rect 124312 114504 124364 114510
rect 124312 114446 124364 114452
rect 124220 114436 124272 114442
rect 124220 114378 124272 114384
rect 125612 68626 125640 170614
rect 126256 117298 126284 253234
rect 126348 202162 126376 254526
rect 126980 253972 127032 253978
rect 126980 253914 127032 253920
rect 126888 253292 126940 253298
rect 126888 253234 126940 253240
rect 126900 253026 126928 253234
rect 126888 253020 126940 253026
rect 126888 252962 126940 252968
rect 126704 251456 126756 251462
rect 126704 251398 126756 251404
rect 126612 251252 126664 251258
rect 126612 251194 126664 251200
rect 126428 248600 126480 248606
rect 126428 248542 126480 248548
rect 126440 203590 126468 248542
rect 126520 248464 126572 248470
rect 126520 248406 126572 248412
rect 126532 231130 126560 248406
rect 126624 233918 126652 251194
rect 126716 234802 126744 251398
rect 126704 234796 126756 234802
rect 126704 234738 126756 234744
rect 126612 233912 126664 233918
rect 126612 233854 126664 233860
rect 126520 231124 126572 231130
rect 126520 231066 126572 231072
rect 126428 203584 126480 203590
rect 126428 203526 126480 203532
rect 126336 202156 126388 202162
rect 126336 202098 126388 202104
rect 126336 198212 126388 198218
rect 126336 198154 126388 198160
rect 126348 197538 126376 198154
rect 126336 197532 126388 197538
rect 126336 197474 126388 197480
rect 126244 117292 126296 117298
rect 126244 117234 126296 117240
rect 125520 68598 125640 68626
rect 123760 67380 123812 67386
rect 123760 67322 123812 67328
rect 123668 66156 123720 66162
rect 123668 66098 123720 66104
rect 125520 66094 125548 68598
rect 125324 66088 125376 66094
rect 125324 66030 125376 66036
rect 125508 66088 125560 66094
rect 125508 66030 125560 66036
rect 123484 65884 123536 65890
rect 123484 65826 123536 65832
rect 124128 65884 124180 65890
rect 124128 65826 124180 65832
rect 111156 65816 111208 65822
rect 111156 65758 111208 65764
rect 121460 65816 121512 65822
rect 121460 65758 121512 65764
rect 122104 65816 122156 65822
rect 122104 65758 122156 65764
rect 124140 65686 124168 65826
rect 124128 65680 124180 65686
rect 124128 65622 124180 65628
rect 125336 65278 125364 66030
rect 126348 65754 126376 197474
rect 126888 170672 126940 170678
rect 126888 170614 126940 170620
rect 126900 169930 126928 170614
rect 126888 169924 126940 169930
rect 126888 169866 126940 169872
rect 126796 117292 126848 117298
rect 126796 117234 126848 117240
rect 126808 116686 126836 117234
rect 126796 116680 126848 116686
rect 126796 116622 126848 116628
rect 126992 114306 127020 253914
rect 133328 253224 133380 253230
rect 133328 253166 133380 253172
rect 130384 251864 130436 251870
rect 130384 251806 130436 251812
rect 127808 251660 127860 251666
rect 127808 251602 127860 251608
rect 127716 250164 127768 250170
rect 127716 250106 127768 250112
rect 127624 247784 127676 247790
rect 127624 247726 127676 247732
rect 127636 247246 127664 247726
rect 127624 247240 127676 247246
rect 127624 247182 127676 247188
rect 127072 198416 127124 198422
rect 127072 198358 127124 198364
rect 127084 197402 127112 198358
rect 127072 197396 127124 197402
rect 127072 197338 127124 197344
rect 127636 114374 127664 247182
rect 127728 201482 127756 250106
rect 127820 237590 127848 251602
rect 129740 250572 129792 250578
rect 129740 250514 129792 250520
rect 129752 250034 129780 250514
rect 129740 250028 129792 250034
rect 129740 249970 129792 249976
rect 129004 245744 129056 245750
rect 129004 245686 129056 245692
rect 127808 237584 127860 237590
rect 127808 237526 127860 237532
rect 129016 236774 129044 245686
rect 130396 236842 130424 251806
rect 131118 251288 131174 251297
rect 131118 251223 131120 251232
rect 131172 251223 131174 251232
rect 131856 251252 131908 251258
rect 131120 251194 131172 251200
rect 131856 251194 131908 251200
rect 130476 250504 130528 250510
rect 130476 250446 130528 250452
rect 130488 249966 130516 250446
rect 130568 250028 130620 250034
rect 130568 249970 130620 249976
rect 130476 249960 130528 249966
rect 130476 249902 130528 249908
rect 130384 236836 130436 236842
rect 130384 236778 130436 236784
rect 129004 236768 129056 236774
rect 129004 236710 129056 236716
rect 127716 201476 127768 201482
rect 127716 201418 127768 201424
rect 129740 198348 129792 198354
rect 129740 198290 129792 198296
rect 129752 197470 129780 198290
rect 129740 197464 129792 197470
rect 129740 197406 129792 197412
rect 130384 197464 130436 197470
rect 130384 197406 130436 197412
rect 127716 197396 127768 197402
rect 127716 197338 127768 197344
rect 127624 114368 127676 114374
rect 127624 114310 127676 114316
rect 126980 114300 127032 114306
rect 126980 114242 127032 114248
rect 127636 114102 127664 114310
rect 127624 114096 127676 114102
rect 127624 114038 127676 114044
rect 127728 74534 127756 197338
rect 128360 196716 128412 196722
rect 128360 196658 128412 196664
rect 127808 169244 127860 169250
rect 127808 169186 127860 169192
rect 127636 74506 127756 74534
rect 127636 67250 127664 74506
rect 127820 68134 127848 169186
rect 127808 68128 127860 68134
rect 127808 68070 127860 68076
rect 127624 67244 127676 67250
rect 127624 67186 127676 67192
rect 127636 66842 127664 67186
rect 127624 66836 127676 66842
rect 127624 66778 127676 66784
rect 126888 65884 126940 65890
rect 126888 65826 126940 65832
rect 126900 65754 126928 65826
rect 126336 65748 126388 65754
rect 126336 65690 126388 65696
rect 126888 65748 126940 65754
rect 126888 65690 126940 65696
rect 125324 65272 125376 65278
rect 125324 65214 125376 65220
rect 111064 64320 111116 64326
rect 111064 64262 111116 64268
rect 110328 64116 110380 64122
rect 110328 64058 110380 64064
rect 128372 16574 128400 196658
rect 130396 67046 130424 197406
rect 130488 119678 130516 249902
rect 130580 122398 130608 249970
rect 131120 198280 131172 198286
rect 131120 198222 131172 198228
rect 131132 197606 131160 198222
rect 131120 197600 131172 197606
rect 131120 197542 131172 197548
rect 131764 197600 131816 197606
rect 131764 197542 131816 197548
rect 130568 122392 130620 122398
rect 130568 122334 130620 122340
rect 131120 121440 131172 121446
rect 131118 121408 131120 121417
rect 131172 121408 131174 121417
rect 131118 121343 131174 121352
rect 130476 119672 130528 119678
rect 130476 119614 130528 119620
rect 131776 67114 131804 197542
rect 131868 121417 131896 251194
rect 133142 247616 133198 247625
rect 133142 247551 133198 247560
rect 131948 237584 132000 237590
rect 131948 237526 132000 237532
rect 131960 122466 131988 237526
rect 131948 122460 132000 122466
rect 131948 122402 132000 122408
rect 131854 121408 131910 121417
rect 131854 121343 131910 121352
rect 133156 114238 133184 247551
rect 133236 234796 133288 234802
rect 133236 234738 133288 234744
rect 133248 120018 133276 234738
rect 133340 232626 133368 253166
rect 142804 252884 142856 252890
rect 142804 252826 142856 252832
rect 134524 250640 134576 250646
rect 134524 250582 134576 250588
rect 134536 249830 134564 250582
rect 140044 249892 140096 249898
rect 140044 249834 140096 249840
rect 134524 249824 134576 249830
rect 134524 249766 134576 249772
rect 133786 247616 133842 247625
rect 133786 247551 133842 247560
rect 133800 247178 133828 247551
rect 133788 247172 133840 247178
rect 133788 247114 133840 247120
rect 133328 232620 133380 232626
rect 133328 232562 133380 232568
rect 133328 169040 133380 169046
rect 133328 168982 133380 168988
rect 133236 120012 133288 120018
rect 133236 119954 133288 119960
rect 133144 114232 133196 114238
rect 133144 114174 133196 114180
rect 132500 106344 132552 106350
rect 132500 106286 132552 106292
rect 131764 67108 131816 67114
rect 131764 67050 131816 67056
rect 130384 67040 130436 67046
rect 130384 66982 130436 66988
rect 132512 16574 132540 106286
rect 133340 66026 133368 168982
rect 134536 117994 134564 249766
rect 137284 244996 137336 245002
rect 137284 244938 137336 244944
rect 137296 244526 137324 244938
rect 137284 244520 137336 244526
rect 137284 244462 137336 244468
rect 137296 238754 137324 244462
rect 137296 238726 137416 238754
rect 134616 232824 134668 232830
rect 134616 232766 134668 232772
rect 134628 231946 134656 232766
rect 134616 231940 134668 231946
rect 134616 231882 134668 231888
rect 134628 119610 134656 231882
rect 137284 198144 137336 198150
rect 137284 198086 137336 198092
rect 137296 197674 137324 198086
rect 137284 197668 137336 197674
rect 137284 197610 137336 197616
rect 134708 171896 134760 171902
rect 134708 171838 134760 171844
rect 134720 171222 134748 171838
rect 134708 171216 134760 171222
rect 134708 171158 134760 171164
rect 134616 119604 134668 119610
rect 134616 119546 134668 119552
rect 134536 117966 134656 117994
rect 134628 115938 134656 117966
rect 134616 115932 134668 115938
rect 134616 115874 134668 115880
rect 134628 115394 134656 115874
rect 134616 115388 134668 115394
rect 134616 115330 134668 115336
rect 133328 66020 133380 66026
rect 133328 65962 133380 65968
rect 133788 66020 133840 66026
rect 133788 65962 133840 65968
rect 133800 65754 133828 65962
rect 133788 65748 133840 65754
rect 133788 65690 133840 65696
rect 134720 65618 134748 171158
rect 135168 119944 135220 119950
rect 135168 119886 135220 119892
rect 135180 119610 135208 119886
rect 135168 119604 135220 119610
rect 135168 119546 135220 119552
rect 137296 66978 137324 197610
rect 137388 117230 137416 238726
rect 138664 232756 138716 232762
rect 138664 232698 138716 232704
rect 138676 231878 138704 232698
rect 138664 231872 138716 231878
rect 138664 231814 138716 231820
rect 137928 206440 137980 206446
rect 137928 206382 137980 206388
rect 137940 200114 137968 206382
rect 137940 200086 138060 200114
rect 138032 199986 138060 200086
rect 138020 199980 138072 199986
rect 138020 199922 138072 199928
rect 137376 117224 137428 117230
rect 137376 117166 137428 117172
rect 137388 116754 137416 117166
rect 137376 116748 137428 116754
rect 137376 116690 137428 116696
rect 138032 113174 138060 199922
rect 138676 118658 138704 231814
rect 139400 225004 139452 225010
rect 139400 224946 139452 224952
rect 138112 118652 138164 118658
rect 138112 118594 138164 118600
rect 138664 118652 138716 118658
rect 138664 118594 138716 118600
rect 138124 118114 138152 118594
rect 138112 118108 138164 118114
rect 138112 118050 138164 118056
rect 137940 113146 138060 113174
rect 137940 112538 137968 113146
rect 137928 112532 137980 112538
rect 137928 112474 137980 112480
rect 137940 95198 137968 112474
rect 137928 95192 137980 95198
rect 137928 95134 137980 95140
rect 137284 66972 137336 66978
rect 137284 66914 137336 66920
rect 135168 66020 135220 66026
rect 135168 65962 135220 65968
rect 135180 65618 135208 65962
rect 134708 65612 134760 65618
rect 134708 65554 134760 65560
rect 135168 65612 135220 65618
rect 135168 65554 135220 65560
rect 139412 16574 139440 224946
rect 140056 121310 140084 249834
rect 140778 232520 140834 232529
rect 140778 232455 140834 232464
rect 140792 232082 140820 232455
rect 140780 232076 140832 232082
rect 140780 232018 140832 232024
rect 141424 232076 141476 232082
rect 141424 232018 141476 232024
rect 140780 174548 140832 174554
rect 140780 174490 140832 174496
rect 140792 173942 140820 174490
rect 140780 173936 140832 173942
rect 140780 173878 140832 173884
rect 140044 121304 140096 121310
rect 140044 121246 140096 121252
rect 140780 113960 140832 113966
rect 140780 113902 140832 113908
rect 140792 113801 140820 113902
rect 141436 113801 141464 232018
rect 141516 173936 141568 173942
rect 141516 173878 141568 173884
rect 140778 113792 140834 113801
rect 140778 113727 140834 113736
rect 141422 113792 141478 113801
rect 141422 113727 141478 113736
rect 141528 67425 141556 173878
rect 142816 114034 142844 252826
rect 142908 121174 142936 254526
rect 151084 254516 151136 254522
rect 151084 254458 151136 254464
rect 148324 253088 148376 253094
rect 148324 253030 148376 253036
rect 144184 251320 144236 251326
rect 144184 251262 144236 251268
rect 142988 213988 143040 213994
rect 142988 213930 143040 213936
rect 143000 189174 143028 213930
rect 142988 189168 143040 189174
rect 142988 189110 143040 189116
rect 143448 170536 143500 170542
rect 143448 170478 143500 170484
rect 143460 169998 143488 170478
rect 142988 169992 143040 169998
rect 142988 169934 143040 169940
rect 143448 169992 143500 169998
rect 143448 169934 143500 169940
rect 142896 121168 142948 121174
rect 142896 121110 142948 121116
rect 142804 114028 142856 114034
rect 142804 113970 142856 113976
rect 141514 67416 141570 67425
rect 141514 67351 141570 67360
rect 143000 66910 143028 169934
rect 143448 121440 143500 121446
rect 143448 121382 143500 121388
rect 143460 121174 143488 121382
rect 144196 121378 144224 251262
rect 146944 250164 146996 250170
rect 146944 250106 146996 250112
rect 144276 229220 144328 229226
rect 144276 229162 144328 229168
rect 144288 213926 144316 229162
rect 144920 214668 144972 214674
rect 144920 214610 144972 214616
rect 145932 214668 145984 214674
rect 145932 214610 145984 214616
rect 144276 213920 144328 213926
rect 144276 213862 144328 213868
rect 144276 189168 144328 189174
rect 144276 189110 144328 189116
rect 144288 165238 144316 189110
rect 144276 165232 144328 165238
rect 144276 165174 144328 165180
rect 144828 165232 144880 165238
rect 144828 165174 144880 165180
rect 144184 121372 144236 121378
rect 144184 121314 144236 121320
rect 144196 121174 144224 121314
rect 143448 121168 143500 121174
rect 143448 121110 143500 121116
rect 144184 121168 144236 121174
rect 144184 121110 144236 121116
rect 143446 114064 143502 114073
rect 143446 113999 143448 114008
rect 143500 113999 143502 114008
rect 143448 113970 143500 113976
rect 144840 85542 144868 165174
rect 144932 115870 144960 214610
rect 145944 213994 145972 214610
rect 145932 213988 145984 213994
rect 145932 213930 145984 213936
rect 146956 120970 146984 250106
rect 147588 239488 147640 239494
rect 147588 239430 147640 239436
rect 147600 238814 147628 239430
rect 147588 238808 147640 238814
rect 147588 238750 147640 238756
rect 147600 125526 147628 238750
rect 147036 125520 147088 125526
rect 147036 125462 147088 125468
rect 147588 125520 147640 125526
rect 147588 125462 147640 125468
rect 147048 124914 147076 125462
rect 147036 124908 147088 124914
rect 147036 124850 147088 124856
rect 146944 120964 146996 120970
rect 146944 120906 146996 120912
rect 144920 115864 144972 115870
rect 144920 115806 144972 115812
rect 145564 115864 145616 115870
rect 145564 115806 145616 115812
rect 145576 115122 145604 115806
rect 145564 115116 145616 115122
rect 145564 115058 145616 115064
rect 145576 98025 145604 115058
rect 147048 103494 147076 124850
rect 148336 121378 148364 253030
rect 150440 231124 150492 231130
rect 150440 231066 150492 231072
rect 150452 230654 150480 231066
rect 150440 230648 150492 230654
rect 150440 230590 150492 230596
rect 148416 216028 148468 216034
rect 148416 215970 148468 215976
rect 148428 165170 148456 215970
rect 148416 165164 148468 165170
rect 148416 165106 148468 165112
rect 148968 165164 149020 165170
rect 148968 165106 149020 165112
rect 148324 121372 148376 121378
rect 148324 121314 148376 121320
rect 148336 121106 148364 121314
rect 148324 121100 148376 121106
rect 148324 121042 148376 121048
rect 147036 103488 147088 103494
rect 147036 103430 147088 103436
rect 145562 98016 145618 98025
rect 145562 97951 145618 97960
rect 144828 85536 144880 85542
rect 144828 85478 144880 85484
rect 144840 84862 144868 85478
rect 144828 84856 144880 84862
rect 144828 84798 144880 84804
rect 148980 71670 149008 165106
rect 150452 112305 150480 230590
rect 150532 186992 150584 186998
rect 150532 186934 150584 186940
rect 150544 186386 150572 186934
rect 150532 186380 150584 186386
rect 150532 186322 150584 186328
rect 151096 120834 151124 254458
rect 153212 254454 153240 702406
rect 169668 576904 169720 576910
rect 169668 576846 169720 576852
rect 169576 484424 169628 484430
rect 169576 484366 169628 484372
rect 169024 298172 169076 298178
rect 169024 298114 169076 298120
rect 167736 257372 167788 257378
rect 167736 257314 167788 257320
rect 155224 254720 155276 254726
rect 155224 254662 155276 254668
rect 153200 254448 153252 254454
rect 153200 254390 153252 254396
rect 153844 254448 153896 254454
rect 153844 254390 153896 254396
rect 152462 250608 152518 250617
rect 152462 250543 152518 250552
rect 152476 250102 152504 250543
rect 152464 250096 152516 250102
rect 152464 250038 152516 250044
rect 151728 186380 151780 186386
rect 151728 186322 151780 186328
rect 151084 120828 151136 120834
rect 151084 120770 151136 120776
rect 150438 112296 150494 112305
rect 150438 112231 150494 112240
rect 150452 110362 150480 112231
rect 150440 110356 150492 110362
rect 150440 110298 150492 110304
rect 151740 80714 151768 186322
rect 152476 113898 152504 250038
rect 153856 219366 153884 254390
rect 155236 253978 155264 254662
rect 167276 254380 167328 254386
rect 167276 254322 167328 254328
rect 167184 254312 167236 254318
rect 167184 254254 167236 254260
rect 155224 253972 155276 253978
rect 155224 253914 155276 253920
rect 153844 219360 153896 219366
rect 153844 219302 153896 219308
rect 154580 214600 154632 214606
rect 154580 214542 154632 214548
rect 152556 200184 152608 200190
rect 152556 200126 152608 200132
rect 152568 165102 152596 200126
rect 152556 165096 152608 165102
rect 152556 165038 152608 165044
rect 153108 165096 153160 165102
rect 153108 165038 153160 165044
rect 153014 113928 153070 113937
rect 152464 113892 152516 113898
rect 153014 113863 153016 113872
rect 152464 113834 152516 113840
rect 153068 113863 153070 113872
rect 153016 113834 153068 113840
rect 151728 80708 151780 80714
rect 151728 80650 151780 80656
rect 153120 74526 153148 165038
rect 154592 115666 154620 214542
rect 155236 122534 155264 253914
rect 164148 252952 164200 252958
rect 164148 252894 164200 252900
rect 157984 252000 158036 252006
rect 157984 251942 158036 251948
rect 157996 251394 158024 251942
rect 157984 251388 158036 251394
rect 157984 251330 158036 251336
rect 156604 249144 156656 249150
rect 156604 249086 156656 249092
rect 156616 248674 156644 249086
rect 156604 248668 156656 248674
rect 156604 248610 156656 248616
rect 155684 214600 155736 214606
rect 155684 214542 155736 214548
rect 155696 214062 155724 214542
rect 155684 214056 155736 214062
rect 155684 213998 155736 214004
rect 155868 189780 155920 189786
rect 155868 189722 155920 189728
rect 155880 189174 155908 189722
rect 155868 189168 155920 189174
rect 155868 189110 155920 189116
rect 155224 122528 155276 122534
rect 155224 122470 155276 122476
rect 155236 122262 155264 122470
rect 155224 122256 155276 122262
rect 155224 122198 155276 122204
rect 154580 115660 154632 115666
rect 154580 115602 154632 115608
rect 155224 115660 155276 115666
rect 155224 115602 155276 115608
rect 154592 115054 154620 115602
rect 154580 115048 154632 115054
rect 154580 114990 154632 114996
rect 155236 100570 155264 115602
rect 155224 100564 155276 100570
rect 155224 100506 155276 100512
rect 155880 83502 155908 189110
rect 156616 121038 156644 248610
rect 156788 212560 156840 212566
rect 156788 212502 156840 212508
rect 156696 169108 156748 169114
rect 156696 169050 156748 169056
rect 156708 168434 156736 169050
rect 156696 168428 156748 168434
rect 156696 168370 156748 168376
rect 156604 121032 156656 121038
rect 156604 120974 156656 120980
rect 155868 83496 155920 83502
rect 155868 83438 155920 83444
rect 153108 74520 153160 74526
rect 153108 74462 153160 74468
rect 153120 73953 153148 74462
rect 153106 73944 153162 73953
rect 153106 73879 153162 73888
rect 148968 71664 149020 71670
rect 148968 71606 149020 71612
rect 142988 66904 143040 66910
rect 142988 66846 143040 66852
rect 155880 65482 155908 83438
rect 156708 68542 156736 168370
rect 156800 165617 156828 212502
rect 157340 199572 157392 199578
rect 157340 199514 157392 199520
rect 157352 198150 157380 199514
rect 157340 198144 157392 198150
rect 157340 198086 157392 198092
rect 156880 183592 156932 183598
rect 156880 183534 156932 183540
rect 156892 167414 156920 183534
rect 156880 167408 156932 167414
rect 156880 167350 156932 167356
rect 156786 165608 156842 165617
rect 156786 165543 156842 165552
rect 156800 161474 156828 165543
rect 156800 161446 157288 161474
rect 157260 84182 157288 161446
rect 157996 118590 158024 251330
rect 159364 249076 159416 249082
rect 159364 249018 159416 249024
rect 159376 248606 159404 249018
rect 159364 248600 159416 248606
rect 159364 248542 159416 248548
rect 158076 239420 158128 239426
rect 158076 239362 158128 239368
rect 158088 238882 158116 239362
rect 158076 238876 158128 238882
rect 158076 238818 158128 238824
rect 158088 121038 158116 238818
rect 158720 207664 158772 207670
rect 158720 207606 158772 207612
rect 158732 207058 158760 207606
rect 158720 207052 158772 207058
rect 158720 206994 158772 207000
rect 158168 198144 158220 198150
rect 158168 198086 158220 198092
rect 158076 121032 158128 121038
rect 158076 120974 158128 120980
rect 158088 120766 158116 120974
rect 158076 120760 158128 120766
rect 158076 120702 158128 120708
rect 157340 118584 157392 118590
rect 157340 118526 157392 118532
rect 157984 118584 158036 118590
rect 157984 118526 158036 118532
rect 157352 118046 157380 118526
rect 157340 118040 157392 118046
rect 157340 117982 157392 117988
rect 158180 113174 158208 198086
rect 157996 113146 158208 113174
rect 157996 112402 158024 113146
rect 157984 112396 158036 112402
rect 157984 112338 158036 112344
rect 157996 89690 158024 112338
rect 158732 112334 158760 206994
rect 159376 122330 159404 248542
rect 162124 248464 162176 248470
rect 162124 248406 162176 248412
rect 159456 240780 159508 240786
rect 159456 240722 159508 240728
rect 159468 240174 159496 240722
rect 159456 240168 159508 240174
rect 159456 240110 159508 240116
rect 159364 122324 159416 122330
rect 159364 122266 159416 122272
rect 159468 122194 159496 240110
rect 159548 123412 159600 123418
rect 159548 123354 159600 123360
rect 159456 122188 159508 122194
rect 159456 122130 159508 122136
rect 158720 112328 158772 112334
rect 158720 112270 158772 112276
rect 158732 111858 158760 112270
rect 158720 111852 158772 111858
rect 158720 111794 158772 111800
rect 159364 111852 159416 111858
rect 159364 111794 159416 111800
rect 159376 96626 159404 111794
rect 159560 100638 159588 123354
rect 162136 121242 162164 248406
rect 163504 229900 163556 229906
rect 163504 229842 163556 229848
rect 162400 229356 162452 229362
rect 162400 229298 162452 229304
rect 162216 211540 162268 211546
rect 162216 211482 162268 211488
rect 162124 121236 162176 121242
rect 162124 121178 162176 121184
rect 162228 112266 162256 211482
rect 162308 210860 162360 210866
rect 162308 210802 162360 210808
rect 162320 114782 162348 210802
rect 162412 206378 162440 229298
rect 163516 219434 163544 229842
rect 163504 219428 163556 219434
rect 163504 219370 163556 219376
rect 162860 215960 162912 215966
rect 162860 215902 162912 215908
rect 162400 206372 162452 206378
rect 162400 206314 162452 206320
rect 162400 190528 162452 190534
rect 162400 190470 162452 190476
rect 162412 167550 162440 190470
rect 162400 167544 162452 167550
rect 162400 167486 162452 167492
rect 162492 125044 162544 125050
rect 162492 124986 162544 124992
rect 162400 123344 162452 123350
rect 162400 123286 162452 123292
rect 162308 114776 162360 114782
rect 162308 114718 162360 114724
rect 162308 113484 162360 113490
rect 162308 113426 162360 113432
rect 162216 112260 162268 112266
rect 162216 112202 162268 112208
rect 162124 112192 162176 112198
rect 162030 112160 162086 112169
rect 162124 112134 162176 112140
rect 162030 112095 162086 112104
rect 162044 103494 162072 112095
rect 162032 103488 162084 103494
rect 162032 103430 162084 103436
rect 159548 100632 159600 100638
rect 159548 100574 159600 100580
rect 159364 96620 159416 96626
rect 159364 96562 159416 96568
rect 157984 89684 158036 89690
rect 157984 89626 158036 89632
rect 162136 85542 162164 112134
rect 162228 97918 162256 112202
rect 162216 97912 162268 97918
rect 162216 97854 162268 97860
rect 162320 88330 162348 113426
rect 162412 93838 162440 123286
rect 162504 99346 162532 124986
rect 162584 124976 162636 124982
rect 162584 124918 162636 124924
rect 162596 100706 162624 124918
rect 162872 114850 162900 215902
rect 163504 182232 163556 182238
rect 163504 182174 163556 182180
rect 163516 167822 163544 182174
rect 163596 180872 163648 180878
rect 163596 180814 163648 180820
rect 163504 167816 163556 167822
rect 163504 167758 163556 167764
rect 163608 167482 163636 180814
rect 163964 167748 164016 167754
rect 163964 167690 164016 167696
rect 163596 167476 163648 167482
rect 163596 167418 163648 167424
rect 163780 164756 163832 164762
rect 163780 164698 163832 164704
rect 163688 122324 163740 122330
rect 163688 122266 163740 122272
rect 163700 121786 163728 122266
rect 163688 121780 163740 121786
rect 163688 121722 163740 121728
rect 163700 116618 163728 121722
rect 163688 116612 163740 116618
rect 163688 116554 163740 116560
rect 162860 114844 162912 114850
rect 162860 114786 162912 114792
rect 163504 114844 163556 114850
rect 163504 114786 163556 114792
rect 162676 114776 162728 114782
rect 162676 114718 162728 114724
rect 162584 100700 162636 100706
rect 162584 100642 162636 100648
rect 162492 99340 162544 99346
rect 162492 99282 162544 99288
rect 162688 96529 162716 114718
rect 162768 112124 162820 112130
rect 162768 112066 162820 112072
rect 162780 102134 162808 112066
rect 162768 102128 162820 102134
rect 162768 102070 162820 102076
rect 163516 100706 163544 114786
rect 163504 100700 163556 100706
rect 163504 100642 163556 100648
rect 162674 96520 162730 96529
rect 162674 96455 162730 96464
rect 162400 93832 162452 93838
rect 162400 93774 162452 93780
rect 162308 88324 162360 88330
rect 162308 88266 162360 88272
rect 162124 85536 162176 85542
rect 162124 85478 162176 85484
rect 157248 84176 157300 84182
rect 157248 84118 157300 84124
rect 157260 83570 157288 84118
rect 157248 83564 157300 83570
rect 157248 83506 157300 83512
rect 162124 82884 162176 82890
rect 162124 82826 162176 82832
rect 156696 68536 156748 68542
rect 156696 68478 156748 68484
rect 162136 66230 162164 82826
rect 162216 77308 162268 77314
rect 162216 77250 162268 77256
rect 162124 66224 162176 66230
rect 162124 66166 162176 66172
rect 162228 65550 162256 77250
rect 162400 76084 162452 76090
rect 162400 76026 162452 76032
rect 162308 76016 162360 76022
rect 162308 75958 162360 75964
rect 162320 65958 162348 75958
rect 162308 65952 162360 65958
rect 162308 65894 162360 65900
rect 162412 65618 162440 76026
rect 162860 75948 162912 75954
rect 162860 75890 162912 75896
rect 162872 71602 162900 75890
rect 162860 71596 162912 71602
rect 162860 71538 162912 71544
rect 163410 68912 163466 68921
rect 163410 68847 163466 68856
rect 163424 67969 163452 68847
rect 163792 68746 163820 164698
rect 163872 164688 163924 164694
rect 163872 164630 163924 164636
rect 163884 68785 163912 164630
rect 163976 69018 164004 167690
rect 164056 167612 164108 167618
rect 164056 167554 164108 167560
rect 163964 69012 164016 69018
rect 163964 68954 164016 68960
rect 164068 68921 164096 167554
rect 164160 122330 164188 252894
rect 165528 252816 165580 252822
rect 165528 252758 165580 252764
rect 165436 229424 165488 229430
rect 165436 229366 165488 229372
rect 164884 226364 164936 226370
rect 164884 226306 164936 226312
rect 164896 198694 164924 226306
rect 165448 225622 165476 229366
rect 165436 225616 165488 225622
rect 165436 225558 165488 225564
rect 164976 202904 165028 202910
rect 164976 202846 165028 202852
rect 164884 198688 164936 198694
rect 164884 198630 164936 198636
rect 164884 189100 164936 189106
rect 164884 189042 164936 189048
rect 164896 168065 164924 189042
rect 164882 168056 164938 168065
rect 164882 167991 164938 168000
rect 164884 165028 164936 165034
rect 164884 164970 164936 164976
rect 164148 122324 164200 122330
rect 164148 122266 164200 122272
rect 164146 122088 164202 122097
rect 164146 122023 164202 122032
rect 164160 118658 164188 122023
rect 164148 118652 164200 118658
rect 164148 118594 164200 118600
rect 164792 118108 164844 118114
rect 164792 118050 164844 118056
rect 164698 112296 164754 112305
rect 164698 112231 164754 112240
rect 164712 111897 164740 112231
rect 164698 111888 164754 111897
rect 164698 111823 164754 111832
rect 164804 107506 164832 118050
rect 164792 107500 164844 107506
rect 164792 107442 164844 107448
rect 164896 86970 164924 164970
rect 164988 163538 165016 202846
rect 165434 169552 165490 169561
rect 165434 169487 165490 169496
rect 164976 163532 165028 163538
rect 164976 163474 165028 163480
rect 164976 124160 165028 124166
rect 164976 124102 165028 124108
rect 164988 123146 165016 124102
rect 165252 123684 165304 123690
rect 165252 123626 165304 123632
rect 165160 123616 165212 123622
rect 165160 123558 165212 123564
rect 165068 123548 165120 123554
rect 165068 123490 165120 123496
rect 164976 123140 165028 123146
rect 164976 123082 165028 123088
rect 164988 115326 165016 123082
rect 164976 115320 165028 115326
rect 164976 115262 165028 115268
rect 164976 113416 165028 113422
rect 164976 113358 165028 113364
rect 164988 91050 165016 113358
rect 165080 106282 165108 123490
rect 165172 118114 165200 123558
rect 165160 118108 165212 118114
rect 165160 118050 165212 118056
rect 165264 117994 165292 123626
rect 165344 118856 165396 118862
rect 165344 118798 165396 118804
rect 165172 117966 165292 117994
rect 165172 110430 165200 117966
rect 165356 115954 165384 118798
rect 165264 115926 165384 115954
rect 165264 111790 165292 115926
rect 165344 113280 165396 113286
rect 165344 113222 165396 113228
rect 165252 111784 165304 111790
rect 165252 111726 165304 111732
rect 165160 110424 165212 110430
rect 165160 110366 165212 110372
rect 165356 106282 165384 113222
rect 165068 106276 165120 106282
rect 165068 106218 165120 106224
rect 165344 106276 165396 106282
rect 165344 106218 165396 106224
rect 164976 91044 165028 91050
rect 164976 90986 165028 90992
rect 165068 90364 165120 90370
rect 165068 90306 165120 90312
rect 164148 86964 164200 86970
rect 164148 86906 164200 86912
rect 164884 86964 164936 86970
rect 164884 86906 164936 86912
rect 164160 85678 164188 86906
rect 164148 85672 164200 85678
rect 164148 85614 164200 85620
rect 164054 68912 164110 68921
rect 164054 68847 164110 68856
rect 163870 68776 163926 68785
rect 163780 68740 163832 68746
rect 163870 68711 163926 68720
rect 163780 68682 163832 68688
rect 163410 67960 163466 67969
rect 163410 67895 163466 67904
rect 162400 65612 162452 65618
rect 162400 65554 162452 65560
rect 162216 65544 162268 65550
rect 162216 65486 162268 65492
rect 164160 65482 164188 85614
rect 164884 84856 164936 84862
rect 164884 84798 164936 84804
rect 164792 73364 164844 73370
rect 164792 73306 164844 73312
rect 164804 70310 164832 73306
rect 164896 71534 164924 84798
rect 164976 78804 165028 78810
rect 164976 78746 165028 78752
rect 164884 71528 164936 71534
rect 164884 71470 164936 71476
rect 164792 70304 164844 70310
rect 164792 70246 164844 70252
rect 164988 69850 165016 78746
rect 165080 69970 165108 90306
rect 165160 78804 165212 78810
rect 165160 78746 165212 78752
rect 165172 70242 165200 78746
rect 165448 74534 165476 169487
rect 165540 124166 165568 252758
rect 166816 232688 166868 232694
rect 166816 232630 166868 232636
rect 166828 232014 166856 232630
rect 166908 232144 166960 232150
rect 166908 232086 166960 232092
rect 166816 232008 166868 232014
rect 166816 231950 166868 231956
rect 166264 229764 166316 229770
rect 166264 229706 166316 229712
rect 166276 204950 166304 229706
rect 166356 229696 166408 229702
rect 166356 229638 166408 229644
rect 166368 211818 166396 229638
rect 166448 229628 166500 229634
rect 166448 229570 166500 229576
rect 166460 217326 166488 229570
rect 166724 229560 166776 229566
rect 166724 229502 166776 229508
rect 166540 229492 166592 229498
rect 166540 229434 166592 229440
rect 166552 220794 166580 229434
rect 166736 224942 166764 229502
rect 166724 224936 166776 224942
rect 166724 224878 166776 224884
rect 166540 220788 166592 220794
rect 166540 220730 166592 220736
rect 166448 217320 166500 217326
rect 166448 217262 166500 217268
rect 166356 211812 166408 211818
rect 166356 211754 166408 211760
rect 166264 204944 166316 204950
rect 166264 204886 166316 204892
rect 166356 197668 166408 197674
rect 166356 197610 166408 197616
rect 166264 197532 166316 197538
rect 166264 197474 166316 197480
rect 166276 168978 166304 197474
rect 166368 169522 166396 197610
rect 166448 197600 166500 197606
rect 166448 197542 166500 197548
rect 166460 169726 166488 197542
rect 166540 194676 166592 194682
rect 166540 194618 166592 194624
rect 166448 169720 166500 169726
rect 166448 169662 166500 169668
rect 166356 169516 166408 169522
rect 166356 169458 166408 169464
rect 166264 168972 166316 168978
rect 166264 168914 166316 168920
rect 166552 167793 166580 194618
rect 166632 176724 166684 176730
rect 166632 176666 166684 176672
rect 166644 168162 166672 176666
rect 166632 168156 166684 168162
rect 166632 168098 166684 168104
rect 166538 167784 166594 167793
rect 166538 167719 166594 167728
rect 166356 164960 166408 164966
rect 166356 164902 166408 164908
rect 166264 164824 166316 164830
rect 166264 164766 166316 164772
rect 165528 124160 165580 124166
rect 165528 124102 165580 124108
rect 165986 122224 166042 122233
rect 165986 122159 166042 122168
rect 166000 115938 166028 122159
rect 166172 120624 166224 120630
rect 166172 120566 166224 120572
rect 166080 120420 166132 120426
rect 166080 120362 166132 120368
rect 165988 115932 166040 115938
rect 165988 115874 166040 115880
rect 166092 114306 166120 120362
rect 166184 114442 166212 120566
rect 166172 114436 166224 114442
rect 166172 114378 166224 114384
rect 166080 114300 166132 114306
rect 166080 114242 166132 114248
rect 165528 113348 165580 113354
rect 165528 113290 165580 113296
rect 165540 107642 165568 113290
rect 165528 107636 165580 107642
rect 165528 107578 165580 107584
rect 165528 97980 165580 97986
rect 165528 97922 165580 97928
rect 165540 96694 165568 97922
rect 165528 96688 165580 96694
rect 165528 96630 165580 96636
rect 165356 74506 165476 74534
rect 165160 70236 165212 70242
rect 165160 70178 165212 70184
rect 165252 70236 165304 70242
rect 165252 70178 165304 70184
rect 165068 69964 165120 69970
rect 165068 69906 165120 69912
rect 165264 69850 165292 70178
rect 164988 69822 165292 69850
rect 165356 67561 165384 74506
rect 165540 73386 165568 96630
rect 166172 79348 166224 79354
rect 166172 79290 166224 79296
rect 165448 73358 165568 73386
rect 165342 67552 165398 67561
rect 165342 67487 165398 67496
rect 165448 66842 165476 73358
rect 165528 73296 165580 73302
rect 165528 73238 165580 73244
rect 165540 69902 165568 73238
rect 166080 70440 166132 70446
rect 166080 70382 166132 70388
rect 165528 69896 165580 69902
rect 165528 69838 165580 69844
rect 165526 67552 165582 67561
rect 165526 67487 165582 67496
rect 165540 67153 165568 67487
rect 165526 67144 165582 67153
rect 165526 67079 165582 67088
rect 165436 66836 165488 66842
rect 165436 66778 165488 66784
rect 155868 65476 155920 65482
rect 155868 65418 155920 65424
rect 164148 65476 164200 65482
rect 164148 65418 164200 65424
rect 155880 65346 155908 65418
rect 155868 65340 155920 65346
rect 155868 65282 155920 65288
rect 164884 65340 164936 65346
rect 164884 65282 164936 65288
rect 164896 46918 164924 65282
rect 166092 64394 166120 70382
rect 166184 68898 166212 79290
rect 166276 78742 166304 164766
rect 166368 97986 166396 164902
rect 166724 162172 166776 162178
rect 166724 162114 166776 162120
rect 166538 121952 166594 121961
rect 166538 121887 166594 121896
rect 166448 120080 166500 120086
rect 166448 120022 166500 120028
rect 166460 119882 166488 120022
rect 166448 119876 166500 119882
rect 166448 119818 166500 119824
rect 166448 118924 166500 118930
rect 166448 118866 166500 118872
rect 166460 111722 166488 118866
rect 166552 117298 166580 121887
rect 166632 119740 166684 119746
rect 166632 119682 166684 119688
rect 166540 117292 166592 117298
rect 166540 117234 166592 117240
rect 166644 114510 166672 119682
rect 166632 114504 166684 114510
rect 166632 114446 166684 114452
rect 166448 111716 166500 111722
rect 166448 111658 166500 111664
rect 166356 97980 166408 97986
rect 166356 97922 166408 97928
rect 166448 95260 166500 95266
rect 166448 95202 166500 95208
rect 166356 94580 166408 94586
rect 166356 94522 166408 94528
rect 166264 78736 166316 78742
rect 166264 78678 166316 78684
rect 166276 69086 166304 78678
rect 166264 69080 166316 69086
rect 166264 69022 166316 69028
rect 166264 68944 166316 68950
rect 166184 68892 166264 68898
rect 166184 68886 166316 68892
rect 166184 68870 166304 68886
rect 166276 68105 166304 68870
rect 166262 68096 166318 68105
rect 166262 68031 166318 68040
rect 166368 67289 166396 94522
rect 166460 69766 166488 95202
rect 166540 94512 166592 94518
rect 166540 94454 166592 94460
rect 166552 69834 166580 94454
rect 166632 89004 166684 89010
rect 166632 88946 166684 88952
rect 166540 69828 166592 69834
rect 166540 69770 166592 69776
rect 166448 69760 166500 69766
rect 166448 69702 166500 69708
rect 166644 69630 166672 88946
rect 166736 79354 166764 162114
rect 166828 122058 166856 231950
rect 166816 122052 166868 122058
rect 166816 121994 166868 122000
rect 166828 117978 166856 121994
rect 166920 119746 166948 232086
rect 167000 229832 167052 229838
rect 167000 229774 167052 229780
rect 167012 229265 167040 229774
rect 166998 229256 167054 229265
rect 166998 229191 167054 229200
rect 166908 119740 166960 119746
rect 166908 119682 166960 119688
rect 166906 119640 166962 119649
rect 166906 119575 166962 119584
rect 166816 117972 166868 117978
rect 166816 117914 166868 117920
rect 166920 115258 166948 119575
rect 167012 118402 167040 229191
rect 167092 229084 167144 229090
rect 167092 229026 167144 229032
rect 167104 227905 167132 229026
rect 167090 227896 167146 227905
rect 167090 227831 167146 227840
rect 167090 225856 167146 225865
rect 167090 225791 167146 225800
rect 167104 225010 167132 225791
rect 167092 225004 167144 225010
rect 167092 224946 167144 224952
rect 167092 224868 167144 224874
rect 167092 224810 167144 224816
rect 167104 224505 167132 224810
rect 167090 224496 167146 224505
rect 167090 224431 167146 224440
rect 167090 223136 167146 223145
rect 167090 223071 167146 223080
rect 167104 222222 167132 223071
rect 167092 222216 167144 222222
rect 167092 222158 167144 222164
rect 167092 219360 167144 219366
rect 167092 219302 167144 219308
rect 167104 219065 167132 219302
rect 167090 219056 167146 219065
rect 167090 218991 167146 219000
rect 167092 218000 167144 218006
rect 167092 217942 167144 217948
rect 167104 217705 167132 217942
rect 167090 217696 167146 217705
rect 167090 217631 167146 217640
rect 167090 216336 167146 216345
rect 167090 216271 167146 216280
rect 167104 215966 167132 216271
rect 167092 215960 167144 215966
rect 167092 215902 167144 215908
rect 167196 215098 167224 254254
rect 167288 229094 167316 254322
rect 167644 254244 167696 254250
rect 167644 254186 167696 254192
rect 167288 229066 167408 229094
rect 167196 215070 167316 215098
rect 167182 214976 167238 214985
rect 167182 214911 167238 214920
rect 167090 214296 167146 214305
rect 167090 214231 167146 214240
rect 167104 213994 167132 214231
rect 167196 214062 167224 214911
rect 167184 214056 167236 214062
rect 167184 213998 167236 214004
rect 167092 213988 167144 213994
rect 167092 213930 167144 213936
rect 167090 211576 167146 211585
rect 167090 211511 167092 211520
rect 167144 211511 167146 211520
rect 167092 211482 167144 211488
rect 167288 210905 167316 215070
rect 167380 211585 167408 229066
rect 167550 227216 167606 227225
rect 167550 227151 167606 227160
rect 167564 226370 167592 227151
rect 167552 226364 167604 226370
rect 167552 226306 167604 226312
rect 167460 221468 167512 221474
rect 167460 221410 167512 221416
rect 167472 221105 167500 221410
rect 167458 221096 167514 221105
rect 167458 221031 167514 221040
rect 167366 211576 167422 211585
rect 167366 211511 167422 211520
rect 167090 210896 167146 210905
rect 167090 210831 167092 210840
rect 167144 210831 167146 210840
rect 167274 210896 167330 210905
rect 167274 210831 167330 210840
rect 167092 210802 167144 210808
rect 167472 209774 167500 221031
rect 167656 212945 167684 254186
rect 167748 254182 167776 257314
rect 167736 254176 167788 254182
rect 167736 254118 167788 254124
rect 167748 219745 167776 254118
rect 167828 252748 167880 252754
rect 167828 252690 167880 252696
rect 167840 222465 167868 252690
rect 168288 242208 168340 242214
rect 168288 242150 168340 242156
rect 168196 231124 168248 231130
rect 168196 231066 168248 231072
rect 167826 222456 167882 222465
rect 167826 222391 167882 222400
rect 167734 219736 167790 219745
rect 167734 219671 167790 219680
rect 167642 212936 167698 212945
rect 167642 212871 167698 212880
rect 167196 209746 167500 209774
rect 167090 208176 167146 208185
rect 167090 208111 167146 208120
rect 167104 207058 167132 208111
rect 167092 207052 167144 207058
rect 167092 206994 167144 207000
rect 167090 206816 167146 206825
rect 167090 206751 167146 206760
rect 167104 206446 167132 206751
rect 167092 206440 167144 206446
rect 167092 206382 167144 206388
rect 167092 206304 167144 206310
rect 167092 206246 167144 206252
rect 167104 206145 167132 206246
rect 167090 206136 167146 206145
rect 167090 206071 167146 206080
rect 167092 201476 167144 201482
rect 167092 201418 167144 201424
rect 167104 201385 167132 201418
rect 167090 201376 167146 201385
rect 167090 201311 167146 201320
rect 167196 201226 167224 209746
rect 167366 206136 167422 206145
rect 167366 206071 167422 206080
rect 167276 203584 167328 203590
rect 167276 203526 167328 203532
rect 167288 203425 167316 203526
rect 167274 203416 167330 203425
rect 167274 203351 167330 203360
rect 167104 201198 167224 201226
rect 167288 201210 167316 203351
rect 167276 201204 167328 201210
rect 167104 118538 167132 201198
rect 167276 201146 167328 201152
rect 167380 201090 167408 206071
rect 167458 202736 167514 202745
rect 167458 202671 167514 202680
rect 167472 202162 167500 202671
rect 167460 202156 167512 202162
rect 167460 202098 167512 202104
rect 167196 201062 167408 201090
rect 167196 118658 167224 201062
rect 167276 201000 167328 201006
rect 167276 200942 167328 200948
rect 167288 123758 167316 200942
rect 167366 200016 167422 200025
rect 167366 199951 167422 199960
rect 167380 199510 167408 199951
rect 167368 199504 167420 199510
rect 167368 199446 167420 199452
rect 167368 198144 167420 198150
rect 167368 198086 167420 198092
rect 167380 197985 167408 198086
rect 167366 197976 167422 197985
rect 167366 197911 167422 197920
rect 167368 196648 167420 196654
rect 167366 196616 167368 196625
rect 167420 196616 167422 196625
rect 167366 196551 167422 196560
rect 167368 192500 167420 192506
rect 167368 192442 167420 192448
rect 167380 191865 167408 192442
rect 167366 191856 167422 191865
rect 167366 191791 167422 191800
rect 167366 189816 167422 189825
rect 167366 189751 167422 189760
rect 167380 189174 167408 189751
rect 167368 189168 167420 189174
rect 167368 189110 167420 189116
rect 167366 186416 167422 186425
rect 167366 186351 167368 186360
rect 167420 186351 167422 186360
rect 167368 186322 167420 186328
rect 167368 185632 167420 185638
rect 167368 185574 167420 185580
rect 167380 185065 167408 185574
rect 167366 185056 167422 185065
rect 167366 184991 167422 185000
rect 167368 184884 167420 184890
rect 167368 184826 167420 184832
rect 167380 183705 167408 184826
rect 167366 183696 167422 183705
rect 167366 183631 167422 183640
rect 167368 183524 167420 183530
rect 167368 183466 167420 183472
rect 167380 182345 167408 183466
rect 167366 182336 167422 182345
rect 167366 182271 167422 182280
rect 167472 180794 167500 202098
rect 167380 180766 167500 180794
rect 167380 128354 167408 180766
rect 167458 180296 167514 180305
rect 167458 180231 167514 180240
rect 167472 180130 167500 180231
rect 167460 180124 167512 180130
rect 167460 180066 167512 180072
rect 167460 177336 167512 177342
rect 167460 177278 167512 177284
rect 167472 176905 167500 177278
rect 167458 176896 167514 176905
rect 167458 176831 167514 176840
rect 167656 132494 167684 212871
rect 168208 209778 168236 231066
rect 168196 209772 168248 209778
rect 168196 209714 168248 209720
rect 168208 209545 168236 209714
rect 168194 209536 168250 209545
rect 168194 209471 168250 209480
rect 168300 206825 168328 242150
rect 168932 239420 168984 239426
rect 168932 239362 168984 239368
rect 168286 206816 168342 206825
rect 168286 206751 168342 206760
rect 168196 199436 168248 199442
rect 168196 199378 168248 199384
rect 168208 195265 168236 199378
rect 168944 198257 168972 239362
rect 169036 199442 169064 298114
rect 169116 236700 169168 236706
rect 169116 236642 169168 236648
rect 169024 199436 169076 199442
rect 169024 199378 169076 199384
rect 168930 198248 168986 198257
rect 168930 198183 168986 198192
rect 168288 198008 168340 198014
rect 168288 197950 168340 197956
rect 168194 195256 168250 195265
rect 168194 195191 168250 195200
rect 168300 193225 168328 197950
rect 169024 196036 169076 196042
rect 169024 195978 169076 195984
rect 168286 193216 168342 193225
rect 168286 193151 168342 193160
rect 168104 191140 168156 191146
rect 168104 191082 168156 191088
rect 168116 190505 168144 191082
rect 168102 190496 168158 190505
rect 168102 190431 168158 190440
rect 168286 185056 168342 185065
rect 168286 184991 168342 185000
rect 168194 180296 168250 180305
rect 168194 180231 168250 180240
rect 168104 175976 168156 175982
rect 168104 175918 168156 175924
rect 168116 175545 168144 175918
rect 168102 175536 168158 175545
rect 168102 175471 168158 175480
rect 168104 172508 168156 172514
rect 168104 172450 168156 172456
rect 168116 172145 168144 172450
rect 168102 172136 168158 172145
rect 168102 172071 168158 172080
rect 168102 170776 168158 170785
rect 168102 170711 168158 170720
rect 168116 170406 168144 170711
rect 168104 170400 168156 170406
rect 168104 170342 168156 170348
rect 167920 170264 167972 170270
rect 167920 170206 167972 170212
rect 167932 167618 167960 170206
rect 168012 169788 168064 169794
rect 168012 169730 168064 169736
rect 167920 167612 167972 167618
rect 167920 167554 167972 167560
rect 167656 132466 167960 132494
rect 167380 128326 167684 128354
rect 167276 123752 167328 123758
rect 167276 123694 167328 123700
rect 167276 119332 167328 119338
rect 167276 119274 167328 119280
rect 167288 118833 167316 119274
rect 167274 118824 167330 118833
rect 167274 118759 167330 118768
rect 167184 118652 167236 118658
rect 167184 118594 167236 118600
rect 167104 118510 167592 118538
rect 167012 118374 167224 118402
rect 167090 118280 167146 118289
rect 167090 118215 167146 118224
rect 166998 117600 167054 117609
rect 166998 117535 167054 117544
rect 167012 117434 167040 117535
rect 167104 117502 167132 118215
rect 167092 117496 167144 117502
rect 167092 117438 167144 117444
rect 167000 117428 167052 117434
rect 167000 117370 167052 117376
rect 166998 115560 167054 115569
rect 166998 115495 167054 115504
rect 166908 115252 166960 115258
rect 166908 115194 166960 115200
rect 167012 114986 167040 115495
rect 167196 115002 167224 118374
rect 167000 114980 167052 114986
rect 167000 114922 167052 114928
rect 167104 114974 167224 115002
rect 167104 114714 167132 114974
rect 167184 114912 167236 114918
rect 167182 114880 167184 114889
rect 167236 114880 167238 114889
rect 167182 114815 167238 114824
rect 167092 114708 167144 114714
rect 167092 114650 167144 114656
rect 166908 113212 166960 113218
rect 166908 113154 166960 113160
rect 166920 112470 166948 113154
rect 166908 112464 166960 112470
rect 166908 112406 166960 112412
rect 166998 112160 167054 112169
rect 166998 112095 167054 112104
rect 167012 112062 167040 112095
rect 167000 112056 167052 112062
rect 167000 111998 167052 112004
rect 166906 111888 166962 111897
rect 166906 111823 166962 111832
rect 166920 93265 166948 111823
rect 167000 110356 167052 110362
rect 167000 110298 167052 110304
rect 167012 110265 167040 110298
rect 166998 110256 167054 110265
rect 166998 110191 167054 110200
rect 167104 109585 167132 114650
rect 167564 114578 167592 118510
rect 167656 116074 167684 128326
rect 167828 123752 167880 123758
rect 167828 123694 167880 123700
rect 167736 118652 167788 118658
rect 167736 118594 167788 118600
rect 167644 116068 167696 116074
rect 167644 116010 167696 116016
rect 167552 114572 167604 114578
rect 167552 114514 167604 114520
rect 167564 113174 167592 114514
rect 167472 113146 167592 113174
rect 167090 109576 167146 109585
rect 167090 109511 167146 109520
rect 167000 107636 167052 107642
rect 167000 107578 167052 107584
rect 167012 107545 167040 107578
rect 166998 107536 167054 107545
rect 166998 107471 167054 107480
rect 166998 106720 167054 106729
rect 166998 106655 167054 106664
rect 167012 106350 167040 106655
rect 167000 106344 167052 106350
rect 167000 106286 167052 106292
rect 167472 104854 167500 113146
rect 167552 108384 167604 108390
rect 167552 108326 167604 108332
rect 167460 104848 167512 104854
rect 167460 104790 167512 104796
rect 167000 103488 167052 103494
rect 166998 103456 167000 103465
rect 167052 103456 167054 103465
rect 166998 103391 167054 103400
rect 167000 102128 167052 102134
rect 166998 102096 167000 102105
rect 167052 102096 167054 102105
rect 166998 102031 167054 102040
rect 167458 100736 167514 100745
rect 167458 100671 167460 100680
rect 167512 100671 167514 100680
rect 167460 100642 167512 100648
rect 167092 100564 167144 100570
rect 167092 100506 167144 100512
rect 167104 100065 167132 100506
rect 167090 100056 167146 100065
rect 167090 99991 167146 100000
rect 167564 98705 167592 108326
rect 167550 98696 167606 98705
rect 167550 98631 167606 98640
rect 167184 97912 167236 97918
rect 167182 97880 167184 97889
rect 167236 97880 167238 97889
rect 167182 97815 167238 97824
rect 167000 95192 167052 95198
rect 167000 95134 167052 95140
rect 167012 94625 167040 95134
rect 166998 94616 167054 94625
rect 166998 94551 167054 94560
rect 166906 93256 166962 93265
rect 166906 93191 166962 93200
rect 167274 92576 167330 92585
rect 167274 92511 167330 92520
rect 166998 89856 167054 89865
rect 166998 89791 167054 89800
rect 167012 89758 167040 89791
rect 167000 89752 167052 89758
rect 167000 89694 167052 89700
rect 167184 89684 167236 89690
rect 167184 89626 167236 89632
rect 166998 89040 167054 89049
rect 166998 88975 167054 88984
rect 167012 88398 167040 88975
rect 167196 88505 167224 89626
rect 167182 88496 167238 88505
rect 167182 88431 167238 88440
rect 167000 88392 167052 88398
rect 167000 88334 167052 88340
rect 167092 88324 167144 88330
rect 167092 88266 167144 88272
rect 167104 87825 167132 88266
rect 167090 87816 167146 87825
rect 167090 87751 167146 87760
rect 166998 85640 167054 85649
rect 166998 85575 167000 85584
rect 167052 85575 167054 85584
rect 167000 85546 167052 85552
rect 167092 85536 167144 85542
rect 167092 85478 167144 85484
rect 167104 84425 167132 85478
rect 167090 84416 167146 84425
rect 167090 84351 167146 84360
rect 166816 83564 166868 83570
rect 166816 83506 166868 83512
rect 166724 79348 166776 79354
rect 166724 79290 166776 79296
rect 166724 75200 166776 75206
rect 166724 75142 166776 75148
rect 166736 69902 166764 75142
rect 166724 69896 166776 69902
rect 166724 69838 166776 69844
rect 166632 69624 166684 69630
rect 166828 69601 166856 83506
rect 167000 83496 167052 83502
rect 167000 83438 167052 83444
rect 167012 83065 167040 83438
rect 166998 83056 167054 83065
rect 166998 82991 167054 83000
rect 166908 82136 166960 82142
rect 166908 82078 166960 82084
rect 166920 69698 166948 82078
rect 166998 81560 167054 81569
rect 166998 81495 167054 81504
rect 167012 81462 167040 81495
rect 167000 81456 167052 81462
rect 167000 81398 167052 81404
rect 167000 80708 167052 80714
rect 167000 80650 167052 80656
rect 167012 80345 167040 80650
rect 166998 80336 167054 80345
rect 167054 80294 167132 80322
rect 166998 80271 167054 80280
rect 166998 78840 167054 78849
rect 166998 78775 167000 78784
rect 167052 78775 167054 78784
rect 167000 78746 167052 78752
rect 167104 78418 167132 80294
rect 167012 78390 167132 78418
rect 166908 69692 166960 69698
rect 166908 69634 166960 69640
rect 166632 69566 166684 69572
rect 166814 69592 166870 69601
rect 166814 69527 166870 69536
rect 166354 67280 166410 67289
rect 166354 67215 166410 67224
rect 167012 64598 167040 78390
rect 167090 74760 167146 74769
rect 167090 74695 167146 74704
rect 167104 74594 167132 74695
rect 167092 74588 167144 74594
rect 167092 74530 167144 74536
rect 167090 74080 167146 74089
rect 167090 74015 167146 74024
rect 167104 73234 167132 74015
rect 167182 73400 167238 73409
rect 167182 73335 167238 73344
rect 167196 73302 167224 73335
rect 167184 73296 167236 73302
rect 167184 73238 167236 73244
rect 167092 73228 167144 73234
rect 167092 73170 167144 73176
rect 167090 72040 167146 72049
rect 167090 71975 167146 71984
rect 167104 71806 167132 71975
rect 167092 71800 167144 71806
rect 167092 71742 167144 71748
rect 167000 64592 167052 64598
rect 167000 64534 167052 64540
rect 166080 64388 166132 64394
rect 166080 64330 166132 64336
rect 166092 63646 166120 64330
rect 166080 63640 166132 63646
rect 166080 63582 166132 63588
rect 167012 62898 167040 64534
rect 167000 62892 167052 62898
rect 167000 62834 167052 62840
rect 164884 46912 164936 46918
rect 164884 46854 164936 46860
rect 167288 28286 167316 92511
rect 167656 91202 167684 116010
rect 167748 116006 167776 118594
rect 167736 116000 167788 116006
rect 167736 115942 167788 115948
rect 167748 93945 167776 115942
rect 167840 114646 167868 123694
rect 167932 117366 167960 132466
rect 167920 117360 167972 117366
rect 167920 117302 167972 117308
rect 167828 114640 167880 114646
rect 167828 114582 167880 114588
rect 167840 103514 167868 114582
rect 167932 108390 167960 117302
rect 167920 108384 167972 108390
rect 167920 108326 167972 108332
rect 167920 106276 167972 106282
rect 167920 106218 167972 106224
rect 167932 105505 167960 106218
rect 167918 105496 167974 105505
rect 167918 105431 167974 105440
rect 167840 103486 167960 103514
rect 167734 93936 167790 93945
rect 167790 93894 167868 93922
rect 167734 93871 167790 93880
rect 167734 91216 167790 91225
rect 167656 91174 167734 91202
rect 167734 91151 167790 91160
rect 167644 91044 167696 91050
rect 167644 90986 167696 90992
rect 167656 90545 167684 90986
rect 167642 90536 167698 90545
rect 167642 90471 167698 90480
rect 167748 84194 167776 91151
rect 167840 89026 167868 93894
rect 167932 92585 167960 103486
rect 167918 92576 167974 92585
rect 167918 92511 167974 92520
rect 167840 88998 167960 89026
rect 167748 84166 167868 84194
rect 167642 79520 167698 79529
rect 167642 79455 167698 79464
rect 167460 71460 167512 71466
rect 167460 71402 167512 71408
rect 167472 70417 167500 71402
rect 167458 70408 167514 70417
rect 167458 70343 167514 70352
rect 167472 64734 167500 70343
rect 167460 64728 167512 64734
rect 167460 64670 167512 64676
rect 167472 63578 167500 64670
rect 167656 64258 167684 79455
rect 167734 78160 167790 78169
rect 167734 78095 167790 78104
rect 167748 64802 167776 78095
rect 167736 64796 167788 64802
rect 167736 64738 167788 64744
rect 167644 64252 167696 64258
rect 167644 64194 167696 64200
rect 167460 63572 167512 63578
rect 167460 63514 167512 63520
rect 167656 39370 167684 64194
rect 167748 42090 167776 64738
rect 167840 61402 167868 84166
rect 167828 61396 167880 61402
rect 167828 61338 167880 61344
rect 167736 42084 167788 42090
rect 167736 42026 167788 42032
rect 167644 39364 167696 39370
rect 167644 39306 167696 39312
rect 167276 28280 167328 28286
rect 167276 28222 167328 28228
rect 128372 16546 128952 16574
rect 132512 16546 133000 16574
rect 139412 16546 139624 16574
rect 107660 4820 107712 4826
rect 107660 4762 107712 4768
rect 69112 3460 69164 3466
rect 69112 3402 69164 3408
rect 572 2848 624 2854
rect 572 2790 624 2796
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 584 480 612 2790
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 132972 480 133000 16546
rect 136456 3460 136508 3466
rect 136456 3402 136508 3408
rect 136468 480 136496 3402
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 167932 13122 167960 88998
rect 168024 71466 168052 169730
rect 168012 71460 168064 71466
rect 168012 71402 168064 71408
rect 168010 71360 168066 71369
rect 168010 71295 168066 71304
rect 168024 70446 168052 71295
rect 168116 70689 168144 170342
rect 168208 76945 168236 180231
rect 168300 79529 168328 184991
rect 168932 173936 168984 173942
rect 168932 173878 168984 173884
rect 168746 173496 168802 173505
rect 168746 173431 168802 173440
rect 168760 173194 168788 173431
rect 168748 173188 168800 173194
rect 168748 173130 168800 173136
rect 168748 172576 168800 172582
rect 168748 172518 168800 172524
rect 168656 170332 168708 170338
rect 168656 170274 168708 170280
rect 168668 167754 168696 170274
rect 168760 167929 168788 172518
rect 168944 168201 168972 173878
rect 169036 169114 169064 195978
rect 169128 173505 169156 236642
rect 169300 230784 169352 230790
rect 169300 230726 169352 230732
rect 169208 230716 169260 230722
rect 169208 230658 169260 230664
rect 169114 173496 169170 173505
rect 169114 173431 169170 173440
rect 169024 169108 169076 169114
rect 169024 169050 169076 169056
rect 168930 168192 168986 168201
rect 168930 168127 168986 168136
rect 168746 167920 168802 167929
rect 168746 167855 168802 167864
rect 168656 167748 168708 167754
rect 168656 167690 168708 167696
rect 169024 126268 169076 126274
rect 169024 126210 169076 126216
rect 168654 121816 168710 121825
rect 168654 121751 168710 121760
rect 168470 120592 168526 120601
rect 168470 120527 168526 120536
rect 168378 120320 168434 120329
rect 168378 120255 168434 120264
rect 168392 114238 168420 120255
rect 168484 114374 168512 120527
rect 168564 120352 168616 120358
rect 168564 120294 168616 120300
rect 168472 114368 168524 114374
rect 168472 114310 168524 114316
rect 168380 114232 168432 114238
rect 168380 114174 168432 114180
rect 168576 113830 168604 120294
rect 168668 117230 168696 121751
rect 168656 117224 168708 117230
rect 168656 117166 168708 117172
rect 168930 116104 168986 116113
rect 168930 116039 168986 116048
rect 168564 113824 168616 113830
rect 168564 113766 168616 113772
rect 168944 108905 168972 116039
rect 168930 108896 168986 108905
rect 168930 108831 168986 108840
rect 169036 104825 169064 126210
rect 169116 119876 169168 119882
rect 169116 119818 169168 119824
rect 169128 119406 169156 119818
rect 169116 119400 169168 119406
rect 169116 119342 169168 119348
rect 169220 118289 169248 230658
rect 169206 118280 169262 118289
rect 169206 118215 169262 118224
rect 169312 117042 169340 230726
rect 169392 230580 169444 230586
rect 169392 230522 169444 230528
rect 169128 117014 169340 117042
rect 169128 116142 169156 117014
rect 169116 116136 169168 116142
rect 169114 116104 169116 116113
rect 169168 116104 169170 116113
rect 169114 116039 169170 116048
rect 169298 114200 169354 114209
rect 169298 114135 169354 114144
rect 169116 113552 169168 113558
rect 169116 113494 169168 113500
rect 169128 106185 169156 113494
rect 169312 113218 169340 114135
rect 169300 113212 169352 113218
rect 169300 113154 169352 113160
rect 169114 106176 169170 106185
rect 169114 106111 169170 106120
rect 169208 104848 169260 104854
rect 169022 104816 169078 104825
rect 169208 104790 169260 104796
rect 169022 104751 169078 104760
rect 169220 104145 169248 104790
rect 169206 104136 169262 104145
rect 169206 104071 169262 104080
rect 169022 100736 169078 100745
rect 169022 100671 169078 100680
rect 168930 97880 168986 97889
rect 168930 97815 168986 97824
rect 168840 96620 168892 96626
rect 168840 96562 168892 96568
rect 168852 95305 168880 96562
rect 168838 95296 168894 95305
rect 168838 95231 168894 95240
rect 168286 79520 168342 79529
rect 168286 79455 168342 79464
rect 168286 77480 168342 77489
rect 168286 77415 168342 77424
rect 168194 76936 168250 76945
rect 168194 76871 168250 76880
rect 168102 70680 168158 70689
rect 168102 70615 168158 70624
rect 168012 70440 168064 70446
rect 168012 70382 168064 70388
rect 168116 64530 168144 70615
rect 168208 64666 168236 76871
rect 168300 64870 168328 77415
rect 168288 64864 168340 64870
rect 168288 64806 168340 64812
rect 168196 64660 168248 64666
rect 168196 64602 168248 64608
rect 168104 64524 168156 64530
rect 168104 64466 168156 64472
rect 168116 64190 168144 64466
rect 168104 64184 168156 64190
rect 168104 64126 168156 64132
rect 168208 60110 168236 64602
rect 168196 60104 168248 60110
rect 168196 60046 168248 60052
rect 168300 50386 168328 64806
rect 168852 64394 168880 95231
rect 168840 64388 168892 64394
rect 168840 64330 168892 64336
rect 168944 64326 168972 97815
rect 168932 64320 168984 64326
rect 168932 64262 168984 64268
rect 169036 62830 169064 100671
rect 169114 98696 169170 98705
rect 169114 98631 169170 98640
rect 169024 62824 169076 62830
rect 169024 62766 169076 62772
rect 169128 55894 169156 98631
rect 169220 57254 169248 104071
rect 169312 64258 169340 113154
rect 169404 112849 169432 230522
rect 169484 230512 169536 230518
rect 169484 230454 169536 230460
rect 169390 112840 169446 112849
rect 169390 112775 169446 112784
rect 169404 111994 169432 112775
rect 169392 111988 169444 111994
rect 169392 111930 169444 111936
rect 169404 111858 169432 111930
rect 169392 111852 169444 111858
rect 169392 111794 169444 111800
rect 169496 110809 169524 230454
rect 169588 190505 169616 484366
rect 169574 190496 169630 190505
rect 169574 190431 169630 190440
rect 169680 179353 169708 576846
rect 169772 198014 169800 702406
rect 188344 700528 188396 700534
rect 188344 700470 188396 700476
rect 184204 700460 184256 700466
rect 184204 700402 184256 700408
rect 182824 700392 182876 700398
rect 182824 700334 182876 700340
rect 173164 510672 173216 510678
rect 173164 510614 173216 510620
rect 169852 418192 169904 418198
rect 169852 418134 169904 418140
rect 169760 198008 169812 198014
rect 169760 197950 169812 197956
rect 169864 189009 169892 418134
rect 169944 311908 169996 311914
rect 169944 311850 169996 311856
rect 169956 194585 169984 311850
rect 170036 256012 170088 256018
rect 170036 255954 170088 255960
rect 170048 254794 170076 255954
rect 170036 254788 170088 254794
rect 170036 254730 170088 254736
rect 170048 248414 170076 254730
rect 170048 248386 170168 248414
rect 170036 230648 170088 230654
rect 170036 230590 170088 230596
rect 169942 194576 169998 194585
rect 169942 194511 169998 194520
rect 170048 190454 170076 230590
rect 170140 205057 170168 248386
rect 172612 247716 172664 247722
rect 172612 247658 172664 247664
rect 171140 244928 171192 244934
rect 171140 244870 171192 244876
rect 171152 230518 171180 244870
rect 171232 233164 171284 233170
rect 171232 233106 171284 233112
rect 171244 230625 171272 233106
rect 171230 230616 171286 230625
rect 171230 230551 171286 230560
rect 171140 230512 171192 230518
rect 171140 230454 171192 230460
rect 170680 230444 170732 230450
rect 170680 230386 170732 230392
rect 170692 229772 170720 230386
rect 171152 229786 171180 230454
rect 171152 229758 171350 229786
rect 172624 229772 172652 247658
rect 173176 230450 173204 510614
rect 180064 404388 180116 404394
rect 180064 404330 180116 404336
rect 173992 254108 174044 254114
rect 173992 254050 174044 254056
rect 173900 246492 173952 246498
rect 173900 246434 173952 246440
rect 173164 230444 173216 230450
rect 173164 230386 173216 230392
rect 173912 229772 173940 246434
rect 174004 231266 174032 254050
rect 179420 254040 179472 254046
rect 179420 253982 179472 253988
rect 177304 251388 177356 251394
rect 177304 251330 177356 251336
rect 175464 246424 175516 246430
rect 175464 246366 175516 246372
rect 173992 231260 174044 231266
rect 173992 231202 174044 231208
rect 175188 231260 175240 231266
rect 175188 231202 175240 231208
rect 174004 230586 174032 231202
rect 173992 230580 174044 230586
rect 173992 230522 174044 230528
rect 175200 229772 175228 231202
rect 175476 229786 175504 246366
rect 177316 240786 177344 251330
rect 178038 250472 178094 250481
rect 178038 250407 178094 250416
rect 177304 240780 177356 240786
rect 177304 240722 177356 240728
rect 177120 236836 177172 236842
rect 177120 236778 177172 236784
rect 175476 229758 175858 229786
rect 177132 229772 177160 236778
rect 178052 229786 178080 250407
rect 179432 230790 179460 253982
rect 180076 233170 180104 404330
rect 181444 253020 181496 253026
rect 181444 252962 181496 252968
rect 180064 233164 180116 233170
rect 180064 233106 180116 233112
rect 179420 230784 179472 230790
rect 179420 230726 179472 230732
rect 179432 229786 179460 230726
rect 180076 229786 180104 233106
rect 181456 232626 181484 252962
rect 182836 249801 182864 700334
rect 183652 253564 183704 253570
rect 183652 253506 183704 253512
rect 182178 249792 182234 249801
rect 182178 249727 182234 249736
rect 182822 249792 182878 249801
rect 182822 249727 182878 249736
rect 182192 248414 182220 249727
rect 182192 248386 182496 248414
rect 181444 232620 181496 232626
rect 181444 232562 181496 232568
rect 181628 232552 181680 232558
rect 181628 232494 181680 232500
rect 178052 229758 178434 229786
rect 179432 229758 179722 229786
rect 180076 229758 180366 229786
rect 181640 229772 181668 232494
rect 182468 230722 182496 248386
rect 183558 233200 183614 233209
rect 183558 233135 183614 233144
rect 182456 230716 182508 230722
rect 182456 230658 182508 230664
rect 182468 229786 182496 230658
rect 183572 230654 183600 233135
rect 183560 230648 183612 230654
rect 183560 230590 183612 230596
rect 183664 229786 183692 253506
rect 184216 233209 184244 700402
rect 186964 700324 187016 700330
rect 186964 700266 187016 700272
rect 186976 248414 187004 700266
rect 188356 249762 188384 700470
rect 192484 670744 192536 670750
rect 192484 670686 192536 670692
rect 190460 250164 190512 250170
rect 190460 250106 190512 250112
rect 187700 249756 187752 249762
rect 187700 249698 187752 249704
rect 188344 249756 188396 249762
rect 188344 249698 188396 249704
rect 186976 248386 187096 248414
rect 187068 248033 187096 248386
rect 187054 248024 187110 248033
rect 187054 247959 187110 247968
rect 186136 236836 186188 236842
rect 186136 236778 186188 236784
rect 186148 233238 186176 236778
rect 186136 233232 186188 233238
rect 184202 233200 184258 233209
rect 186136 233174 186188 233180
rect 184202 233135 184258 233144
rect 184848 230648 184900 230654
rect 184848 230590 184900 230596
rect 182468 229758 182942 229786
rect 183586 229758 183692 229786
rect 184860 229772 184888 230590
rect 186148 229772 186176 233174
rect 187068 229786 187096 247959
rect 187712 229786 187740 249698
rect 190472 233986 190500 250106
rect 192496 248414 192524 670686
rect 195244 324352 195296 324358
rect 195244 324294 195296 324300
rect 194600 254584 194652 254590
rect 194600 254526 194652 254532
rect 193220 252816 193272 252822
rect 193220 252758 193272 252764
rect 193232 248414 193260 252758
rect 192496 248386 192616 248414
rect 193232 248386 193536 248414
rect 190644 238876 190696 238882
rect 190644 238818 190696 238824
rect 190460 233980 190512 233986
rect 190460 233922 190512 233928
rect 189356 232688 189408 232694
rect 189356 232630 189408 232636
rect 187068 229758 187450 229786
rect 187712 229758 188094 229786
rect 189368 229772 189396 232630
rect 190656 229772 190684 238818
rect 191012 233980 191064 233986
rect 191012 233922 191064 233928
rect 191024 229786 191052 233922
rect 192588 232082 192616 248386
rect 192576 232076 192628 232082
rect 192576 232018 192628 232024
rect 191024 229758 191314 229786
rect 192588 229772 192616 232018
rect 193508 229786 193536 248386
rect 194612 233986 194640 254526
rect 194692 252952 194744 252958
rect 194692 252894 194744 252900
rect 194704 248414 194732 252894
rect 194704 248386 194824 248414
rect 194600 233980 194652 233986
rect 194600 233922 194652 233928
rect 194796 229786 194824 248386
rect 195256 236842 195284 324294
rect 201512 265674 201540 702986
rect 203524 456816 203576 456822
rect 203524 456758 203576 456764
rect 201500 265668 201552 265674
rect 201500 265610 201552 265616
rect 195980 254516 196032 254522
rect 195980 254458 196032 254464
rect 195992 248414 196020 254458
rect 198740 253088 198792 253094
rect 198740 253030 198792 253036
rect 195992 248386 196664 248414
rect 195244 236836 195296 236842
rect 195244 236778 195296 236784
rect 195428 233980 195480 233986
rect 195428 233922 195480 233928
rect 195440 229786 195468 233922
rect 196636 229786 196664 248386
rect 198372 232552 198424 232558
rect 198372 232494 198424 232500
rect 198384 230654 198412 232494
rect 198372 230648 198424 230654
rect 198372 230590 198424 230596
rect 193508 229758 193890 229786
rect 194796 229758 195178 229786
rect 195440 229758 195822 229786
rect 196636 229758 197110 229786
rect 198384 229772 198412 230590
rect 198752 229786 198780 253030
rect 203536 251190 203564 456758
rect 211160 253972 211212 253978
rect 211160 253914 211212 253920
rect 204904 253428 204956 253434
rect 204904 253370 204956 253376
rect 203064 251184 203116 251190
rect 203064 251126 203116 251132
rect 203524 251184 203576 251190
rect 203524 251126 203576 251132
rect 203076 250102 203104 251126
rect 203064 250096 203116 250102
rect 203064 250038 203116 250044
rect 201500 249960 201552 249966
rect 201500 249902 201552 249908
rect 201512 248414 201540 249902
rect 201512 248386 201632 248414
rect 200120 247240 200172 247246
rect 200120 247182 200172 247188
rect 200132 229786 200160 247182
rect 198752 229758 199042 229786
rect 200132 229758 200330 229786
rect 201604 229772 201632 248386
rect 202880 237584 202932 237590
rect 202880 237526 202932 237532
rect 202892 229772 202920 237526
rect 203076 229786 203104 250038
rect 204916 232082 204944 253370
rect 211068 251320 211120 251326
rect 211068 251262 211120 251268
rect 211080 251190 211108 251262
rect 211068 251184 211120 251190
rect 211068 251126 211120 251132
rect 205732 250028 205784 250034
rect 205732 249970 205784 249976
rect 205744 248414 205772 249970
rect 210424 249892 210476 249898
rect 210424 249834 210476 249840
rect 205744 248386 206416 248414
rect 205640 244316 205692 244322
rect 205640 244258 205692 244264
rect 205652 242214 205680 244258
rect 205640 242208 205692 242214
rect 205640 242150 205692 242156
rect 204904 232076 204956 232082
rect 204904 232018 204956 232024
rect 204916 229786 204944 232018
rect 206100 231940 206152 231946
rect 206100 231882 206152 231888
rect 203076 229758 203550 229786
rect 204838 229758 204944 229786
rect 206112 229772 206140 231882
rect 206388 229786 206416 248386
rect 208952 240780 209004 240786
rect 208952 240722 209004 240728
rect 207664 240168 207716 240174
rect 207664 240110 207716 240116
rect 207676 229786 207704 240110
rect 208964 229786 208992 240722
rect 210436 233170 210464 249834
rect 211172 248414 211200 253914
rect 215944 249824 215996 249830
rect 215944 249766 215996 249772
rect 212540 248668 212592 248674
rect 212540 248610 212592 248616
rect 211172 248386 211292 248414
rect 210424 233164 210476 233170
rect 210424 233106 210476 233112
rect 210608 231872 210660 231878
rect 210608 231814 210660 231820
rect 206388 229758 206770 229786
rect 207676 229758 208058 229786
rect 208964 229758 209346 229786
rect 210620 229772 210648 231814
rect 211264 229772 211292 248386
rect 212552 229772 212580 248610
rect 213368 247172 213420 247178
rect 213368 247114 213420 247120
rect 213380 233102 213408 247114
rect 215956 233238 215984 249766
rect 218072 244526 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 233884 683188 233936 683194
rect 233884 683130 233936 683136
rect 228364 258120 228416 258126
rect 228364 258062 228416 258068
rect 219440 252884 219492 252890
rect 219440 252826 219492 252832
rect 218152 248600 218204 248606
rect 218152 248542 218204 248548
rect 218060 244520 218112 244526
rect 218060 244462 218112 244468
rect 218072 233986 218100 244462
rect 218060 233980 218112 233986
rect 218060 233922 218112 233928
rect 215944 233232 215996 233238
rect 215944 233174 215996 233180
rect 217048 233232 217100 233238
rect 217048 233174 217100 233180
rect 214472 233164 214524 233170
rect 214472 233106 214524 233112
rect 213368 233096 213420 233102
rect 213368 233038 213420 233044
rect 213380 229786 213408 233038
rect 213380 229758 213854 229786
rect 214484 229772 214512 233106
rect 215760 232144 215812 232150
rect 215760 232086 215812 232092
rect 215772 229772 215800 232086
rect 217060 229772 217088 233174
rect 218164 229786 218192 248542
rect 219452 248414 219480 252826
rect 222844 251252 222896 251258
rect 222844 251194 222896 251200
rect 219452 248386 219848 248414
rect 218612 233980 218664 233986
rect 218612 233922 218664 233928
rect 218624 229786 218652 233922
rect 219820 229786 219848 248386
rect 222856 233170 222884 251194
rect 228376 251190 228404 258062
rect 227720 251184 227772 251190
rect 227720 251126 227772 251132
rect 228364 251184 228416 251190
rect 228364 251126 228416 251132
rect 223580 248464 223632 248470
rect 223632 248412 224448 248414
rect 223580 248406 224448 248412
rect 223592 248386 224448 248406
rect 222844 233164 222896 233170
rect 222844 233106 222896 233112
rect 221556 232008 221608 232014
rect 221556 231950 221608 231956
rect 223488 232008 223540 232014
rect 223488 231950 223540 231956
rect 218164 229758 218362 229786
rect 218624 229758 219006 229786
rect 219820 229758 220294 229786
rect 221568 229772 221596 231950
rect 222200 231872 222252 231878
rect 222200 231814 222252 231820
rect 222212 229772 222240 231814
rect 223500 229772 223528 231950
rect 224420 229786 224448 248386
rect 226708 234796 226760 234802
rect 226708 234738 226760 234744
rect 226064 233164 226116 233170
rect 226064 233106 226116 233112
rect 226076 232558 226104 233106
rect 226064 232552 226116 232558
rect 226064 232494 226116 232500
rect 224420 229758 224802 229786
rect 226076 229772 226104 232494
rect 226720 229772 226748 234738
rect 227732 229786 227760 251126
rect 230296 247104 230348 247110
rect 230296 247046 230348 247052
rect 229468 246356 229520 246362
rect 229468 246298 229520 246304
rect 229284 233912 229336 233918
rect 229284 233854 229336 233860
rect 229100 230920 229152 230926
rect 229100 230862 229152 230868
rect 227732 229758 228022 229786
rect 229112 219434 229140 230862
rect 229296 229786 229324 233854
rect 229296 229772 229416 229786
rect 229310 229758 229416 229772
rect 229388 229158 229416 229758
rect 229284 229152 229336 229158
rect 229284 229094 229336 229100
rect 229376 229152 229428 229158
rect 229376 229094 229428 229100
rect 229204 229066 229324 229094
rect 229204 227746 229232 229066
rect 229480 228857 229508 246298
rect 230204 245676 230256 245682
rect 230204 245618 230256 245624
rect 230112 243024 230164 243030
rect 230112 242966 230164 242972
rect 230020 241596 230072 241602
rect 230020 241538 230072 241544
rect 229560 234728 229612 234734
rect 229560 234670 229612 234676
rect 229282 228848 229338 228857
rect 229466 228848 229522 228857
rect 229338 228806 229416 228834
rect 229282 228783 229338 228792
rect 229282 227760 229338 227769
rect 229204 227718 229282 227746
rect 229282 227695 229338 227704
rect 229112 219406 229324 219434
rect 229296 209273 229324 219406
rect 229282 209264 229338 209273
rect 229282 209199 229338 209208
rect 170126 205048 170182 205057
rect 170126 204983 170182 204992
rect 229388 203017 229416 228806
rect 229466 228783 229522 228792
rect 229572 212537 229600 234670
rect 229928 230444 229980 230450
rect 229928 230386 229980 230392
rect 229940 229772 229968 230386
rect 229834 228984 229890 228993
rect 229834 228919 229890 228928
rect 229650 226672 229706 226681
rect 229650 226607 229706 226616
rect 229664 226370 229692 226607
rect 229652 226364 229704 226370
rect 229652 226306 229704 226312
rect 229558 212528 229614 212537
rect 229558 212463 229614 212472
rect 229374 203008 229430 203017
rect 229374 202943 229430 202952
rect 170312 198076 170364 198082
rect 170312 198018 170364 198024
rect 170048 190426 170168 190454
rect 169850 189000 169906 189009
rect 169850 188935 169906 188944
rect 169666 179344 169722 179353
rect 169666 179279 169722 179288
rect 169852 171216 169904 171222
rect 169852 171158 169904 171164
rect 169576 171148 169628 171154
rect 169576 171090 169628 171096
rect 169588 168230 169616 171090
rect 169864 170610 169892 171158
rect 169852 170604 169904 170610
rect 169852 170546 169904 170552
rect 169680 170462 170062 170490
rect 169680 169794 169708 170462
rect 169852 170400 169904 170406
rect 169852 170342 169904 170348
rect 169668 169788 169720 169794
rect 169668 169730 169720 169736
rect 169576 168224 169628 168230
rect 169576 168166 169628 168172
rect 169864 168094 169892 170342
rect 170036 170060 170088 170066
rect 170036 170002 170088 170008
rect 169852 168088 169904 168094
rect 169852 168030 169904 168036
rect 170048 167890 170076 170002
rect 170036 167884 170088 167890
rect 170036 167826 170088 167832
rect 170140 161474 170168 190426
rect 170324 173058 170352 198018
rect 170404 197464 170456 197470
rect 170404 197406 170456 197412
rect 170312 173052 170364 173058
rect 170312 172994 170364 173000
rect 170416 172938 170444 197406
rect 170496 197396 170548 197402
rect 170496 197338 170548 197344
rect 170232 172910 170444 172938
rect 170232 169318 170260 172910
rect 170312 172848 170364 172854
rect 170312 172790 170364 172796
rect 170324 169697 170352 172790
rect 170404 171828 170456 171834
rect 170404 171770 170456 171776
rect 170416 170762 170444 171770
rect 170508 170882 170536 197338
rect 229374 196208 229430 196217
rect 229374 196143 229430 196152
rect 170496 170876 170548 170882
rect 170496 170818 170548 170824
rect 170416 170734 170706 170762
rect 170496 170672 170548 170678
rect 170496 170614 170548 170620
rect 170404 170196 170456 170202
rect 170404 170138 170456 170144
rect 170310 169688 170366 169697
rect 170310 169623 170366 169632
rect 170220 169312 170272 169318
rect 170220 169254 170272 169260
rect 170416 168026 170444 170138
rect 170508 169386 170536 170614
rect 171980 170270 172008 170748
rect 173268 170338 173296 170748
rect 173256 170332 173308 170338
rect 173256 170274 173308 170280
rect 173912 170270 173940 170748
rect 175200 170270 175228 170748
rect 176488 170270 176516 170748
rect 177776 170270 177804 170748
rect 178420 170270 178448 170748
rect 179708 170270 179736 170748
rect 180996 170270 181024 170748
rect 181640 170270 181668 170748
rect 182928 170270 182956 170748
rect 184216 170270 184244 170748
rect 185504 170270 185532 170748
rect 186148 170270 186176 170748
rect 187436 170270 187464 170748
rect 188724 170270 188752 170748
rect 189368 170270 189396 170748
rect 190656 170270 190684 170748
rect 191944 170270 191972 170748
rect 193232 170270 193260 170748
rect 193876 170270 193904 170748
rect 195164 170270 195192 170748
rect 196452 170270 196480 170748
rect 197096 170270 197124 170748
rect 198384 170270 198412 170748
rect 199672 170270 199700 170748
rect 200960 170270 200988 170748
rect 201604 170270 201632 170748
rect 202892 170270 202920 170748
rect 204180 170270 204208 170748
rect 204824 170270 204852 170748
rect 206112 170270 206140 170748
rect 207400 170270 207428 170748
rect 208688 170270 208716 170748
rect 209332 170270 209360 170748
rect 210620 170270 210648 170748
rect 211908 170270 211936 170748
rect 212552 170270 212580 170748
rect 213840 170270 213868 170748
rect 215128 170270 215156 170748
rect 216416 170270 216444 170748
rect 217060 170270 217088 170748
rect 218348 170270 218376 170748
rect 219636 170270 219664 170748
rect 220280 170270 220308 170748
rect 221568 170270 221596 170748
rect 222856 170270 222884 170748
rect 224144 170270 224172 170748
rect 224788 170270 224816 170748
rect 226076 170270 226104 170748
rect 227364 170270 227392 170748
rect 228824 170400 228876 170406
rect 228666 170326 228772 170354
rect 228824 170342 228876 170348
rect 171968 170264 172020 170270
rect 171968 170206 172020 170212
rect 173900 170264 173952 170270
rect 173900 170206 173952 170212
rect 175188 170264 175240 170270
rect 175188 170206 175240 170212
rect 176476 170264 176528 170270
rect 176476 170206 176528 170212
rect 177764 170264 177816 170270
rect 177764 170206 177816 170212
rect 178408 170264 178460 170270
rect 178408 170206 178460 170212
rect 179696 170264 179748 170270
rect 179696 170206 179748 170212
rect 180984 170264 181036 170270
rect 180984 170206 181036 170212
rect 181628 170264 181680 170270
rect 181628 170206 181680 170212
rect 182916 170264 182968 170270
rect 182916 170206 182968 170212
rect 184204 170264 184256 170270
rect 184204 170206 184256 170212
rect 185492 170264 185544 170270
rect 185492 170206 185544 170212
rect 186136 170264 186188 170270
rect 186136 170206 186188 170212
rect 187424 170264 187476 170270
rect 187424 170206 187476 170212
rect 188712 170264 188764 170270
rect 188712 170206 188764 170212
rect 189356 170264 189408 170270
rect 189356 170206 189408 170212
rect 190644 170264 190696 170270
rect 190644 170206 190696 170212
rect 191932 170264 191984 170270
rect 191932 170206 191984 170212
rect 193220 170264 193272 170270
rect 193220 170206 193272 170212
rect 193864 170264 193916 170270
rect 193864 170206 193916 170212
rect 195152 170264 195204 170270
rect 195152 170206 195204 170212
rect 196440 170264 196492 170270
rect 196440 170206 196492 170212
rect 197084 170264 197136 170270
rect 197084 170206 197136 170212
rect 198372 170264 198424 170270
rect 198372 170206 198424 170212
rect 199660 170264 199712 170270
rect 199660 170206 199712 170212
rect 200948 170264 201000 170270
rect 200948 170206 201000 170212
rect 201592 170264 201644 170270
rect 201592 170206 201644 170212
rect 202880 170264 202932 170270
rect 202880 170206 202932 170212
rect 204168 170264 204220 170270
rect 204168 170206 204220 170212
rect 204812 170264 204864 170270
rect 204812 170206 204864 170212
rect 206100 170264 206152 170270
rect 206100 170206 206152 170212
rect 207388 170264 207440 170270
rect 207388 170206 207440 170212
rect 208676 170264 208728 170270
rect 208676 170206 208728 170212
rect 209320 170264 209372 170270
rect 209320 170206 209372 170212
rect 210608 170264 210660 170270
rect 210608 170206 210660 170212
rect 211896 170264 211948 170270
rect 211896 170206 211948 170212
rect 212540 170264 212592 170270
rect 212540 170206 212592 170212
rect 213828 170264 213880 170270
rect 213828 170206 213880 170212
rect 215116 170264 215168 170270
rect 215116 170206 215168 170212
rect 216404 170264 216456 170270
rect 216404 170206 216456 170212
rect 217048 170264 217100 170270
rect 217048 170206 217100 170212
rect 218336 170264 218388 170270
rect 218336 170206 218388 170212
rect 219624 170264 219676 170270
rect 219624 170206 219676 170212
rect 220268 170264 220320 170270
rect 220268 170206 220320 170212
rect 221556 170264 221608 170270
rect 221556 170206 221608 170212
rect 222844 170264 222896 170270
rect 222844 170206 222896 170212
rect 224132 170264 224184 170270
rect 224132 170206 224184 170212
rect 224776 170264 224828 170270
rect 224776 170206 224828 170212
rect 226064 170264 226116 170270
rect 226064 170206 226116 170212
rect 227352 170264 227404 170270
rect 227352 170206 227404 170212
rect 173900 169992 173952 169998
rect 173900 169934 173952 169940
rect 175188 169992 175240 169998
rect 175188 169934 175240 169940
rect 175280 169992 175332 169998
rect 175280 169934 175332 169940
rect 177764 169992 177816 169998
rect 177764 169934 177816 169940
rect 178408 169992 178460 169998
rect 178408 169934 178460 169940
rect 179696 169992 179748 169998
rect 179696 169934 179748 169940
rect 180984 169992 181036 169998
rect 180984 169934 181036 169940
rect 181628 169992 181680 169998
rect 181628 169934 181680 169940
rect 182916 169992 182968 169998
rect 182916 169934 182968 169940
rect 184204 169992 184256 169998
rect 184204 169934 184256 169940
rect 185492 169992 185544 169998
rect 185492 169934 185544 169940
rect 186136 169992 186188 169998
rect 186136 169934 186188 169940
rect 187424 169992 187476 169998
rect 187424 169934 187476 169940
rect 188712 169992 188764 169998
rect 188712 169934 188764 169940
rect 189356 169992 189408 169998
rect 189356 169934 189408 169940
rect 189448 169992 189500 169998
rect 189448 169934 189500 169940
rect 191932 169992 191984 169998
rect 191932 169934 191984 169940
rect 193220 169992 193272 169998
rect 193220 169934 193272 169940
rect 193864 169992 193916 169998
rect 193864 169934 193916 169940
rect 195152 169992 195204 169998
rect 195152 169934 195204 169940
rect 196440 169992 196492 169998
rect 196440 169934 196492 169940
rect 196532 169992 196584 169998
rect 196532 169934 196584 169940
rect 198372 169992 198424 169998
rect 198372 169934 198424 169940
rect 199660 169992 199712 169998
rect 199660 169934 199712 169940
rect 201408 169992 201460 169998
rect 201408 169934 201460 169940
rect 201592 169992 201644 169998
rect 201592 169934 201644 169940
rect 202880 169992 202932 169998
rect 202880 169934 202932 169940
rect 204168 169992 204220 169998
rect 204168 169934 204220 169940
rect 204812 169992 204864 169998
rect 204812 169934 204864 169940
rect 206100 169992 206152 169998
rect 206100 169934 206152 169940
rect 207388 169992 207440 169998
rect 207388 169934 207440 169940
rect 208676 169992 208728 169998
rect 208676 169934 208728 169940
rect 210608 169992 210660 169998
rect 210608 169934 210660 169940
rect 211896 169992 211948 169998
rect 211896 169934 211948 169940
rect 212540 169992 212592 169998
rect 212540 169934 212592 169940
rect 213828 169992 213880 169998
rect 213828 169934 213880 169940
rect 215116 169992 215168 169998
rect 215116 169934 215168 169940
rect 216404 169992 216456 169998
rect 216404 169934 216456 169940
rect 217048 169992 217100 169998
rect 217048 169934 217100 169940
rect 218336 169992 218388 169998
rect 218336 169934 218388 169940
rect 219624 169992 219676 169998
rect 219624 169934 219676 169940
rect 220268 169992 220320 169998
rect 220268 169934 220320 169940
rect 221556 169992 221608 169998
rect 221556 169934 221608 169940
rect 222844 169992 222896 169998
rect 222844 169934 222896 169940
rect 224776 169992 224828 169998
rect 224776 169934 224828 169940
rect 226064 169992 226116 169998
rect 226064 169934 226116 169940
rect 227352 169992 227404 169998
rect 227352 169934 227404 169940
rect 170956 169924 171008 169930
rect 170956 169866 171008 169872
rect 170496 169380 170548 169386
rect 170496 169322 170548 169328
rect 170968 168337 170996 169866
rect 171048 169856 171100 169862
rect 171048 169798 171100 169804
rect 171060 168366 171088 169798
rect 173912 169590 173940 169934
rect 175200 169590 175228 169934
rect 173900 169584 173952 169590
rect 173900 169526 173952 169532
rect 175188 169584 175240 169590
rect 175188 169526 175240 169532
rect 175200 169017 175228 169526
rect 175186 169008 175242 169017
rect 175186 168943 175242 168952
rect 175292 168366 175320 169934
rect 171048 168360 171100 168366
rect 170954 168328 171010 168337
rect 171048 168302 171100 168308
rect 175280 168360 175332 168366
rect 175280 168302 175332 168308
rect 170954 168263 171010 168272
rect 170404 168020 170456 168026
rect 170404 167962 170456 167968
rect 177776 167686 177804 169934
rect 178420 168910 178448 169934
rect 178408 168904 178460 168910
rect 178408 168846 178460 168852
rect 177764 167680 177816 167686
rect 177764 167622 177816 167628
rect 179708 167482 179736 169934
rect 179696 167476 179748 167482
rect 179696 167418 179748 167424
rect 180996 164762 181024 169934
rect 181168 169448 181220 169454
rect 181168 169390 181220 169396
rect 181180 167958 181208 169390
rect 181168 167952 181220 167958
rect 181168 167894 181220 167900
rect 180984 164756 181036 164762
rect 180984 164698 181036 164704
rect 181640 164694 181668 169934
rect 182928 167929 182956 169934
rect 182914 167920 182970 167929
rect 182914 167855 182970 167864
rect 182928 167346 182956 167855
rect 182916 167340 182968 167346
rect 182916 167282 182968 167288
rect 184216 164830 184244 169934
rect 184940 168904 184992 168910
rect 184940 168846 184992 168852
rect 184952 168337 184980 168846
rect 184938 168328 184994 168337
rect 184938 168263 184994 168272
rect 185504 167414 185532 169934
rect 186148 168910 186176 169934
rect 186136 168904 186188 168910
rect 186136 168846 186188 168852
rect 187436 168434 187464 169934
rect 187424 168428 187476 168434
rect 187424 168370 187476 168376
rect 185492 167408 185544 167414
rect 185492 167350 185544 167356
rect 188724 165034 188752 169934
rect 189368 167618 189396 169934
rect 189460 169182 189488 169934
rect 189448 169176 189500 169182
rect 189448 169118 189500 169124
rect 189356 167612 189408 167618
rect 189356 167554 189408 167560
rect 188712 165028 188764 165034
rect 188712 164970 188764 164976
rect 184204 164824 184256 164830
rect 184204 164766 184256 164772
rect 181628 164688 181680 164694
rect 181628 164630 181680 164636
rect 191944 162178 191972 169934
rect 193232 168065 193260 169934
rect 193218 168056 193274 168065
rect 193218 167991 193274 168000
rect 193232 167482 193260 167991
rect 193220 167476 193272 167482
rect 193220 167418 193272 167424
rect 193876 164966 193904 169934
rect 195164 167822 195192 169934
rect 196452 168366 196480 169934
rect 196544 169250 196572 169934
rect 198384 169561 198412 169934
rect 198370 169552 198426 169561
rect 198370 169487 198426 169496
rect 198384 169454 198412 169487
rect 198372 169448 198424 169454
rect 198372 169390 198424 169396
rect 196532 169244 196584 169250
rect 196532 169186 196584 169192
rect 196440 168360 196492 168366
rect 199672 168337 199700 169934
rect 201420 168978 201448 169934
rect 201408 168972 201460 168978
rect 201408 168914 201460 168920
rect 196440 168302 196492 168308
rect 199658 168328 199714 168337
rect 199658 168263 199714 168272
rect 195152 167816 195204 167822
rect 195152 167758 195204 167764
rect 195244 167748 195296 167754
rect 195244 167690 195296 167696
rect 193864 164960 193916 164966
rect 193864 164902 193916 164908
rect 191932 162172 191984 162178
rect 191932 162114 191984 162120
rect 170048 161446 170168 161474
rect 170048 132494 170076 161446
rect 170048 132466 170168 132494
rect 170140 128354 170168 132466
rect 170048 128326 170168 128354
rect 169668 127628 169720 127634
rect 169668 127570 169720 127576
rect 169680 126274 169708 127570
rect 169668 126268 169720 126274
rect 169668 126210 169720 126216
rect 169760 121712 169812 121718
rect 169760 121654 169812 121660
rect 169942 121680 169998 121689
rect 169772 120850 169800 121654
rect 169942 121615 169998 121624
rect 169852 121508 169904 121514
rect 169852 121450 169904 121456
rect 169588 120822 169800 120850
rect 169588 119218 169616 120822
rect 169760 120692 169812 120698
rect 169760 120634 169812 120640
rect 169772 120170 169800 120634
rect 169680 120142 169800 120170
rect 169680 119746 169708 120142
rect 169864 120034 169892 121450
rect 169956 120290 169984 121615
rect 169944 120284 169996 120290
rect 169944 120226 169996 120232
rect 169772 120006 169892 120034
rect 169772 119950 169800 120006
rect 169760 119944 169812 119950
rect 169760 119886 169812 119892
rect 169852 119944 169904 119950
rect 169852 119886 169904 119892
rect 169864 119746 169892 119886
rect 169668 119740 169720 119746
rect 169668 119682 169720 119688
rect 169852 119740 169904 119746
rect 169852 119682 169904 119688
rect 170048 119626 170076 128326
rect 183560 126268 183612 126274
rect 183560 126210 183612 126216
rect 174544 124228 174596 124234
rect 174544 124170 174596 124176
rect 170956 122664 171008 122670
rect 170956 122606 171008 122612
rect 170968 120086 170996 122606
rect 173256 122324 173308 122330
rect 173256 122266 173308 122272
rect 173268 121038 173296 122266
rect 173256 121032 173308 121038
rect 173256 120974 173308 120980
rect 170956 120080 171008 120086
rect 170956 120022 171008 120028
rect 171968 119944 172020 119950
rect 171060 119882 171364 119898
rect 171968 119886 172020 119892
rect 171048 119876 171364 119882
rect 171100 119870 171364 119876
rect 171048 119818 171100 119824
rect 171336 119748 171364 119870
rect 171980 119748 172008 119886
rect 172440 119882 172652 119898
rect 172428 119876 172652 119882
rect 172480 119870 172652 119876
rect 172428 119818 172480 119824
rect 172624 119748 172652 119870
rect 173268 119748 173296 120974
rect 174556 120970 174584 124170
rect 183572 124166 183600 126210
rect 182916 124160 182968 124166
rect 182916 124102 182968 124108
rect 183560 124160 183612 124166
rect 183560 124102 183612 124108
rect 175832 123140 175884 123146
rect 175832 123082 175884 123088
rect 175280 121780 175332 121786
rect 175280 121722 175332 121728
rect 174544 120964 174596 120970
rect 174544 120906 174596 120912
rect 174556 119748 174584 120906
rect 175292 120290 175320 121722
rect 175280 120284 175332 120290
rect 175280 120226 175332 120232
rect 175186 120184 175242 120193
rect 175186 120119 175242 120128
rect 175200 119748 175228 120119
rect 175844 119748 175872 123082
rect 179696 122596 179748 122602
rect 179696 122538 179748 122544
rect 178406 121952 178462 121961
rect 178406 121887 178462 121896
rect 177120 121440 177172 121446
rect 177120 121382 177172 121388
rect 177132 120494 177160 121382
rect 177764 120828 177816 120834
rect 177764 120770 177816 120776
rect 177120 120488 177172 120494
rect 177120 120430 177172 120436
rect 176476 120284 176528 120290
rect 176476 120226 176528 120232
rect 176488 119748 176516 120226
rect 177132 119748 177160 120430
rect 177776 119748 177804 120770
rect 178420 119748 178448 121887
rect 179708 121378 179736 122538
rect 181812 122460 181864 122466
rect 181812 122402 181864 122408
rect 181824 121854 181852 122402
rect 181812 121848 181864 121854
rect 181812 121790 181864 121796
rect 180982 121680 181038 121689
rect 180982 121615 181038 121624
rect 179696 121372 179748 121378
rect 179696 121314 179748 121320
rect 179708 119748 179736 121314
rect 180338 120592 180394 120601
rect 180338 120527 180394 120536
rect 180352 119748 180380 120527
rect 180996 119748 181024 121615
rect 181824 121258 181852 121790
rect 181640 121230 181852 121258
rect 181640 119748 181668 121230
rect 182270 120456 182326 120465
rect 182270 120391 182326 120400
rect 182284 119748 182312 120391
rect 182928 120222 182956 124102
rect 195256 122834 195284 167690
rect 195336 167680 195388 167686
rect 195336 167622 195388 167628
rect 195072 122806 195284 122834
rect 187700 122596 187752 122602
rect 187700 122538 187752 122544
rect 187424 122528 187476 122534
rect 187424 122470 187476 122476
rect 184756 122392 184808 122398
rect 184756 122334 184808 122340
rect 184768 121990 184796 122334
rect 185492 122188 185544 122194
rect 185492 122130 185544 122136
rect 184756 121984 184808 121990
rect 184756 121926 184808 121932
rect 183560 121508 183612 121514
rect 183560 121450 183612 121456
rect 182916 120216 182968 120222
rect 182916 120158 182968 120164
rect 182928 119748 182956 120158
rect 183572 119748 183600 121450
rect 184768 120578 184796 121926
rect 184848 121712 184900 121718
rect 184848 121654 184900 121660
rect 184860 120698 184888 121654
rect 184848 120692 184900 120698
rect 184848 120634 184900 120640
rect 184768 120550 184888 120578
rect 184860 119748 184888 120550
rect 185504 120222 185532 122130
rect 186778 122088 186834 122097
rect 186778 122023 186834 122032
rect 186136 121780 186188 121786
rect 186136 121722 186188 121728
rect 185492 120216 185544 120222
rect 185492 120158 185544 120164
rect 185504 119748 185532 120158
rect 186148 119748 186176 121722
rect 186228 121576 186280 121582
rect 186228 121518 186280 121524
rect 186240 121106 186268 121518
rect 186320 121508 186372 121514
rect 186320 121450 186372 121456
rect 186332 121242 186360 121450
rect 186320 121236 186372 121242
rect 186320 121178 186372 121184
rect 186228 121100 186280 121106
rect 186228 121042 186280 121048
rect 186792 120562 186820 122023
rect 187436 121922 187464 122470
rect 187424 121916 187476 121922
rect 187424 121858 187476 121864
rect 186780 120556 186832 120562
rect 186780 120498 186832 120504
rect 186792 119748 186820 120498
rect 187436 119748 187464 121858
rect 187712 120834 187740 122538
rect 191932 122256 191984 122262
rect 191286 122224 191342 122233
rect 188068 122188 188120 122194
rect 191932 122198 191984 122204
rect 191286 122159 191342 122168
rect 188068 122130 188120 122136
rect 188080 121582 188108 122130
rect 190644 121712 190696 121718
rect 190644 121654 190696 121660
rect 188068 121576 188120 121582
rect 188068 121518 188120 121524
rect 187700 120828 187752 120834
rect 187700 120770 187752 120776
rect 188080 119748 188108 121518
rect 190000 121304 190052 121310
rect 190000 121246 190052 121252
rect 188710 120320 188766 120329
rect 188710 120255 188766 120264
rect 188724 119748 188752 120255
rect 190012 119748 190040 121246
rect 190656 119748 190684 121654
rect 191300 119748 191328 122159
rect 191944 119748 191972 122198
rect 193864 122052 193916 122058
rect 193864 121994 193916 122000
rect 192574 121816 192630 121825
rect 192574 121751 192630 121760
rect 192588 119748 192616 121751
rect 193128 121508 193180 121514
rect 193128 121450 193180 121456
rect 193140 121417 193168 121450
rect 193126 121408 193182 121417
rect 193126 121343 193182 121352
rect 193218 120728 193274 120737
rect 193218 120663 193274 120672
rect 193232 120154 193260 120663
rect 193876 120358 193904 121994
rect 195072 120426 195100 122806
rect 195348 120986 195376 167622
rect 201420 162178 201448 168914
rect 201604 167890 201632 169934
rect 202892 168162 202920 169934
rect 203432 168360 203484 168366
rect 203432 168302 203484 168308
rect 202880 168156 202932 168162
rect 202880 168098 202932 168104
rect 201592 167884 201644 167890
rect 201592 167826 201644 167832
rect 202236 166320 202288 166326
rect 202236 166262 202288 166268
rect 202144 164960 202196 164966
rect 202144 164902 202196 164908
rect 201500 163532 201552 163538
rect 201500 163474 201552 163480
rect 201408 162172 201460 162178
rect 201408 162114 201460 162120
rect 199936 160744 199988 160750
rect 199936 160686 199988 160692
rect 199948 122834 199976 160686
rect 200488 124976 200540 124982
rect 200488 124918 200540 124924
rect 200028 124840 200080 124846
rect 200028 124782 200080 124788
rect 199856 122806 199976 122834
rect 197728 122664 197780 122670
rect 197728 122606 197780 122612
rect 196440 121780 196492 121786
rect 196440 121722 196492 121728
rect 196452 121582 196480 121722
rect 196440 121576 196492 121582
rect 196440 121518 196492 121524
rect 195164 120958 195376 120986
rect 195164 120630 195192 120958
rect 195152 120624 195204 120630
rect 195152 120566 195204 120572
rect 195060 120420 195112 120426
rect 195060 120362 195112 120368
rect 193864 120352 193916 120358
rect 193864 120294 193916 120300
rect 193220 120148 193272 120154
rect 193220 120090 193272 120096
rect 193232 119748 193260 120090
rect 193876 119748 193904 120294
rect 195164 119748 195192 120566
rect 195796 120420 195848 120426
rect 195796 120362 195848 120368
rect 195808 119748 195836 120362
rect 196452 119748 196480 121518
rect 197084 121508 197136 121514
rect 197084 121450 197136 121456
rect 197096 119748 197124 121450
rect 197740 119898 197768 122606
rect 198832 122188 198884 122194
rect 198832 122130 198884 122136
rect 198372 121168 198424 121174
rect 198372 121110 198424 121116
rect 197740 119882 197860 119898
rect 197740 119876 197872 119882
rect 197740 119870 197820 119876
rect 197740 119748 197768 119870
rect 197820 119818 197872 119824
rect 198384 119748 198412 121110
rect 198844 119882 198872 122130
rect 199856 121650 199884 122806
rect 199016 121644 199068 121650
rect 199016 121586 199068 121592
rect 199844 121644 199896 121650
rect 199844 121586 199896 121592
rect 198832 119876 198884 119882
rect 198832 119818 198884 119824
rect 199028 119748 199056 121586
rect 199660 119944 199712 119950
rect 199660 119886 199712 119892
rect 199672 119748 199700 119886
rect 169680 119612 170076 119626
rect 169680 119598 170062 119612
rect 169680 119338 169708 119598
rect 170678 119368 170734 119377
rect 169668 119332 169720 119338
rect 170678 119303 170734 119312
rect 169668 119274 169720 119280
rect 169588 119190 169800 119218
rect 169772 118590 169800 119190
rect 169760 118584 169812 118590
rect 169760 118526 169812 118532
rect 169574 116104 169630 116113
rect 169574 116039 169630 116048
rect 169482 110800 169538 110809
rect 169482 110735 169538 110744
rect 169496 110498 169524 110735
rect 169484 110492 169536 110498
rect 169484 110434 169536 110440
rect 169390 109576 169446 109585
rect 169390 109511 169446 109520
rect 169300 64252 169352 64258
rect 169300 64194 169352 64200
rect 169404 61470 169432 109511
rect 169482 100056 169538 100065
rect 169482 99991 169538 100000
rect 169392 61464 169444 61470
rect 169392 61406 169444 61412
rect 169208 57248 169260 57254
rect 169208 57190 169260 57196
rect 169116 55888 169168 55894
rect 169116 55830 169168 55836
rect 168288 50380 168340 50386
rect 168288 50322 168340 50328
rect 169496 49026 169524 99991
rect 169588 62966 169616 116039
rect 200040 113098 200068 124782
rect 200396 124772 200448 124778
rect 200396 124714 200448 124720
rect 200304 124636 200356 124642
rect 200304 124578 200356 124584
rect 200212 123276 200264 123282
rect 200212 123218 200264 123224
rect 200118 119368 200174 119377
rect 200118 119303 200174 119312
rect 200132 118862 200160 119303
rect 200120 118856 200172 118862
rect 200120 118798 200172 118804
rect 200224 113218 200252 123218
rect 200316 113286 200344 124578
rect 200304 113280 200356 113286
rect 200304 113222 200356 113228
rect 200212 113212 200264 113218
rect 200212 113154 200264 113160
rect 200118 113112 200174 113121
rect 200040 113070 200118 113098
rect 200118 113047 200174 113056
rect 200302 113112 200358 113121
rect 200302 113047 200358 113056
rect 200316 112962 200344 113047
rect 200040 112934 200344 112962
rect 169668 111852 169720 111858
rect 169668 111794 169720 111800
rect 169576 62960 169628 62966
rect 169576 62902 169628 62908
rect 169484 49020 169536 49026
rect 169484 48962 169536 48968
rect 169680 15910 169708 111794
rect 169850 106176 169906 106185
rect 169850 106111 169906 106120
rect 169758 88496 169814 88505
rect 169758 88431 169814 88440
rect 169772 24138 169800 88431
rect 169864 61538 169892 106111
rect 200040 86034 200068 112934
rect 200120 112872 200172 112878
rect 200120 112814 200172 112820
rect 200212 112872 200264 112878
rect 200212 112814 200264 112820
rect 200132 104417 200160 112814
rect 200118 104408 200174 104417
rect 200118 104343 200174 104352
rect 200118 98288 200174 98297
rect 200118 98223 200174 98232
rect 200132 86154 200160 98223
rect 200224 95577 200252 112814
rect 200408 110537 200436 124714
rect 200394 110528 200450 110537
rect 200394 110463 200450 110472
rect 200500 109002 200528 124918
rect 200948 121984 201000 121990
rect 200948 121926 201000 121932
rect 200764 121848 200816 121854
rect 200764 121790 200816 121796
rect 200580 119944 200632 119950
rect 200580 119886 200632 119892
rect 200592 118998 200620 119886
rect 200580 118992 200632 118998
rect 200580 118934 200632 118940
rect 200304 108996 200356 109002
rect 200304 108938 200356 108944
rect 200488 108996 200540 109002
rect 200488 108938 200540 108944
rect 200316 108497 200344 108938
rect 200302 108488 200358 108497
rect 200302 108423 200358 108432
rect 200776 104174 200804 121790
rect 200960 113830 200988 121926
rect 200948 113824 201000 113830
rect 200948 113766 201000 113772
rect 200764 104168 200816 104174
rect 200764 104110 200816 104116
rect 200210 95568 200266 95577
rect 200210 95503 200266 95512
rect 201406 95568 201462 95577
rect 201406 95503 201462 95512
rect 201420 95266 201448 95503
rect 201408 95260 201460 95266
rect 201408 95202 201460 95208
rect 200210 94888 200266 94897
rect 200210 94823 200266 94832
rect 200224 86170 200252 94823
rect 200302 92848 200358 92857
rect 200302 92783 200358 92792
rect 200316 89714 200344 92783
rect 200316 89686 200436 89714
rect 200120 86148 200172 86154
rect 200224 86142 200344 86170
rect 200120 86090 200172 86096
rect 200118 86048 200174 86057
rect 200040 86006 200118 86034
rect 200118 85983 200174 85992
rect 200118 85640 200174 85649
rect 200040 85598 200118 85626
rect 198832 70712 198884 70718
rect 198738 70680 198794 70689
rect 198096 70644 198148 70650
rect 198832 70654 198884 70660
rect 198738 70615 198794 70624
rect 198096 70586 198148 70592
rect 170034 70408 170090 70417
rect 170034 70343 170090 70352
rect 198108 70258 198136 70586
rect 170692 68066 170720 70244
rect 171336 68921 171364 70244
rect 171796 70230 171994 70258
rect 172638 70230 173020 70258
rect 171796 69018 171824 70230
rect 171784 69012 171836 69018
rect 171784 68954 171836 68960
rect 171322 68912 171378 68921
rect 171322 68847 171378 68856
rect 170496 68060 170548 68066
rect 170496 68002 170548 68008
rect 170680 68060 170732 68066
rect 170680 68002 170732 68008
rect 170404 63640 170456 63646
rect 170404 63582 170456 63588
rect 169944 63572 169996 63578
rect 169944 63514 169996 63520
rect 169852 61532 169904 61538
rect 169852 61474 169904 61480
rect 169956 60042 169984 63514
rect 169944 60036 169996 60042
rect 169944 59978 169996 59984
rect 170416 44878 170444 63582
rect 170508 55962 170536 68002
rect 170496 55956 170548 55962
rect 170496 55898 170548 55904
rect 170404 44872 170456 44878
rect 170404 44814 170456 44820
rect 171796 33794 171824 68954
rect 171874 68912 171930 68921
rect 171874 68847 171930 68856
rect 171888 47598 171916 68847
rect 172992 68406 173020 70230
rect 172980 68400 173032 68406
rect 172980 68342 173032 68348
rect 172992 64874 173020 68342
rect 173268 66065 173296 70244
rect 173912 67182 173940 70244
rect 174556 68241 174584 70244
rect 174542 68232 174598 68241
rect 174542 68167 174598 68176
rect 173900 67176 173952 67182
rect 173900 67118 173952 67124
rect 173254 66056 173310 66065
rect 173254 65991 173310 66000
rect 172992 64846 173204 64874
rect 171876 47592 171928 47598
rect 171876 47534 171928 47540
rect 171784 33788 171836 33794
rect 171784 33730 171836 33736
rect 169760 24132 169812 24138
rect 169760 24074 169812 24080
rect 169668 15904 169720 15910
rect 169668 15846 169720 15852
rect 173176 14482 173204 64846
rect 173164 14476 173216 14482
rect 173164 14418 173216 14424
rect 167920 13116 167972 13122
rect 167920 13058 167972 13064
rect 174556 4826 174584 68167
rect 175844 67454 175872 70244
rect 175936 70230 176502 70258
rect 177146 70230 177436 70258
rect 175936 68338 175964 70230
rect 177302 68776 177358 68785
rect 177408 68746 177436 70230
rect 177776 68785 177804 70244
rect 178040 69080 178092 69086
rect 178040 69022 178092 69028
rect 177762 68776 177818 68785
rect 177302 68711 177358 68720
rect 177396 68740 177448 68746
rect 175924 68332 175976 68338
rect 175924 68274 175976 68280
rect 175832 67448 175884 67454
rect 175832 67390 175884 67396
rect 175844 65414 175872 67390
rect 175832 65408 175884 65414
rect 175832 65350 175884 65356
rect 175936 11762 175964 68274
rect 175924 11756 175976 11762
rect 175924 11698 175976 11704
rect 174544 4820 174596 4826
rect 174544 4762 174596 4768
rect 177316 3466 177344 68711
rect 177762 68711 177818 68720
rect 177396 68682 177448 68688
rect 177408 3670 177436 68682
rect 178052 49094 178080 69022
rect 178420 65929 178448 70244
rect 179064 69086 179092 70244
rect 179052 69080 179104 69086
rect 179052 69022 179104 69028
rect 179708 68377 179736 70244
rect 179694 68368 179750 68377
rect 179694 68303 179750 68312
rect 180062 68368 180118 68377
rect 180062 68303 180118 68312
rect 178406 65920 178462 65929
rect 178406 65855 178462 65864
rect 178040 49088 178092 49094
rect 178040 49030 178092 49036
rect 180076 4962 180104 68303
rect 180996 66774 181024 70244
rect 181456 70230 181654 70258
rect 182298 70230 182680 70258
rect 181456 68542 181484 70230
rect 181444 68536 181496 68542
rect 181444 68478 181496 68484
rect 180984 66768 181036 66774
rect 180984 66710 181036 66716
rect 180064 4956 180116 4962
rect 180064 4898 180116 4904
rect 181456 4894 181484 68478
rect 182652 65482 182680 70230
rect 182928 67318 182956 70244
rect 182916 67312 182968 67318
rect 182916 67254 182968 67260
rect 183572 65822 183600 70244
rect 184216 68950 184244 70244
rect 184204 68944 184256 68950
rect 184204 68886 184256 68892
rect 183560 65816 183612 65822
rect 183560 65758 183612 65764
rect 182640 65476 182692 65482
rect 182640 65418 182692 65424
rect 182652 64874 182680 65418
rect 182652 64846 182864 64874
rect 182836 6866 182864 64846
rect 182824 6860 182876 6866
rect 182824 6802 182876 6808
rect 181444 4888 181496 4894
rect 181444 4830 181496 4836
rect 177396 3664 177448 3670
rect 177396 3606 177448 3612
rect 184216 3534 184244 68886
rect 184860 65686 184888 70244
rect 185596 70230 186162 70258
rect 186806 70230 187004 70258
rect 185596 66842 185624 70230
rect 186976 68270 187004 70230
rect 187436 68474 187464 70244
rect 188094 70230 188384 70258
rect 187424 68468 187476 68474
rect 187424 68410 187476 68416
rect 186964 68264 187016 68270
rect 186964 68206 187016 68212
rect 185584 66836 185636 66842
rect 185584 66778 185636 66784
rect 184848 65680 184900 65686
rect 184848 65622 184900 65628
rect 185596 7682 185624 66778
rect 186976 46238 187004 68206
rect 187436 67182 187464 68410
rect 188356 68202 188384 70230
rect 188344 68196 188396 68202
rect 188344 68138 188396 68144
rect 187424 67176 187476 67182
rect 187424 67118 187476 67124
rect 187436 64874 187464 67118
rect 187436 64846 187648 64874
rect 186964 46232 187016 46238
rect 186964 46174 187016 46180
rect 185584 7676 185636 7682
rect 185584 7618 185636 7624
rect 187620 5030 187648 64846
rect 188356 18630 188384 68138
rect 188724 67561 188752 70244
rect 189092 70230 189382 70258
rect 189092 68921 189120 70230
rect 189078 68912 189134 68921
rect 189078 68847 189134 68856
rect 189092 68513 189120 68847
rect 189078 68504 189134 68513
rect 189078 68439 189134 68448
rect 188710 67552 188766 67561
rect 188710 67487 188766 67496
rect 190012 65890 190040 70244
rect 190366 68912 190422 68921
rect 190366 68847 190422 68856
rect 190000 65884 190052 65890
rect 190000 65826 190052 65832
rect 190380 31074 190408 68847
rect 191300 66094 191328 70244
rect 191944 66162 191972 70244
rect 192588 68950 192616 70244
rect 192576 68944 192628 68950
rect 192576 68886 192628 68892
rect 192588 68649 192616 68886
rect 193232 68814 193260 70244
rect 193220 68808 193272 68814
rect 193220 68750 193272 68756
rect 192574 68640 192630 68649
rect 192574 68575 192630 68584
rect 193232 68542 193260 68750
rect 193876 68678 193904 70244
rect 193864 68672 193916 68678
rect 193864 68614 193916 68620
rect 194416 68672 194468 68678
rect 194416 68614 194468 68620
rect 193220 68536 193272 68542
rect 193220 68478 193272 68484
rect 194324 68536 194376 68542
rect 194324 68478 194376 68484
rect 191932 66156 191984 66162
rect 191932 66098 191984 66104
rect 191104 66088 191156 66094
rect 191104 66030 191156 66036
rect 191288 66088 191340 66094
rect 191288 66030 191340 66036
rect 191116 33114 191144 66030
rect 194336 64874 194364 68478
rect 194428 66858 194456 68614
rect 194520 67046 194548 70244
rect 194508 67040 194560 67046
rect 194508 66982 194560 66988
rect 194428 66830 194548 66858
rect 194336 64846 194456 64874
rect 194428 51746 194456 64846
rect 194416 51740 194468 51746
rect 194416 51682 194468 51688
rect 194520 37942 194548 66830
rect 195164 65754 195192 70244
rect 195244 69896 195296 69902
rect 195296 69844 195468 69850
rect 195244 69838 195468 69844
rect 195256 69834 195468 69838
rect 195256 69828 195480 69834
rect 195256 69822 195428 69828
rect 195428 69770 195480 69776
rect 196452 67114 196480 70244
rect 196636 70230 197110 70258
rect 197754 70244 198136 70258
rect 197740 70230 198136 70244
rect 196636 69018 196664 70230
rect 196624 69012 196676 69018
rect 196624 68954 196676 68960
rect 196440 67108 196492 67114
rect 196440 67050 196492 67056
rect 195152 65748 195204 65754
rect 195152 65690 195204 65696
rect 196636 64122 196664 68954
rect 197740 68814 197768 70230
rect 197728 68808 197780 68814
rect 197728 68750 197780 68756
rect 198384 68746 198412 70244
rect 198648 68808 198700 68814
rect 198648 68750 198700 68756
rect 198372 68740 198424 68746
rect 198372 68682 198424 68688
rect 196624 64116 196676 64122
rect 196624 64058 196676 64064
rect 196636 58682 196664 64058
rect 196624 58676 196676 58682
rect 196624 58618 196676 58624
rect 194508 37936 194560 37942
rect 194508 37878 194560 37884
rect 191104 33108 191156 33114
rect 191104 33050 191156 33056
rect 190368 31068 190420 31074
rect 190368 31010 190420 31016
rect 198660 21418 198688 68750
rect 198752 66910 198780 70615
rect 198844 68542 198872 70654
rect 198832 68536 198884 68542
rect 198832 68478 198884 68484
rect 199028 67250 199056 70244
rect 199382 69864 199438 69873
rect 199382 69799 199438 69808
rect 199396 67522 199424 69799
rect 199384 67516 199436 67522
rect 199384 67458 199436 67464
rect 199016 67244 199068 67250
rect 199016 67186 199068 67192
rect 199672 66978 199700 70244
rect 200040 70106 200068 85598
rect 200118 85575 200174 85584
rect 200120 85536 200172 85542
rect 200120 85478 200172 85484
rect 200132 70378 200160 85478
rect 200316 80054 200344 86142
rect 200224 80026 200344 80054
rect 200224 72026 200252 80026
rect 200224 71998 200344 72026
rect 200210 71904 200266 71913
rect 200210 71839 200266 71848
rect 200120 70372 200172 70378
rect 200120 70314 200172 70320
rect 200028 70100 200080 70106
rect 200028 70042 200080 70048
rect 200224 67425 200252 71839
rect 200316 71738 200344 71998
rect 200304 71732 200356 71738
rect 200304 71674 200356 71680
rect 200408 71670 200436 89686
rect 201512 82929 201540 163474
rect 201592 130416 201644 130422
rect 201592 130358 201644 130364
rect 201604 105777 201632 130358
rect 202052 124908 202104 124914
rect 202052 124850 202104 124856
rect 201776 124704 201828 124710
rect 201776 124646 201828 124652
rect 201684 124500 201736 124506
rect 201684 124442 201736 124448
rect 201590 105768 201646 105777
rect 201590 105703 201646 105712
rect 201696 103057 201724 124442
rect 201788 105097 201816 124646
rect 201868 124364 201920 124370
rect 201868 124306 201920 124312
rect 201880 111897 201908 124306
rect 201960 123684 202012 123690
rect 201960 123626 202012 123632
rect 201972 118697 202000 123626
rect 201958 118688 202014 118697
rect 201958 118623 202014 118632
rect 201958 118008 202014 118017
rect 201958 117943 201960 117952
rect 202012 117943 202014 117952
rect 201960 117914 202012 117920
rect 201958 115288 202014 115297
rect 201958 115223 201960 115232
rect 202012 115223 202014 115232
rect 201960 115194 202012 115200
rect 201866 111888 201922 111897
rect 201866 111823 201922 111832
rect 202064 111217 202092 124850
rect 202156 124166 202184 164902
rect 202248 130422 202276 166262
rect 202328 142860 202380 142866
rect 202328 142802 202380 142808
rect 202236 130416 202288 130422
rect 202236 130358 202288 130364
rect 202236 125044 202288 125050
rect 202236 124986 202288 124992
rect 202144 124160 202196 124166
rect 202144 124102 202196 124108
rect 202142 117328 202198 117337
rect 202142 117263 202198 117272
rect 202156 116618 202184 117263
rect 202144 116612 202196 116618
rect 202144 116554 202196 116560
rect 202248 113150 202276 124986
rect 202340 123554 202368 142802
rect 202880 124568 202932 124574
rect 202880 124510 202932 124516
rect 202420 124160 202472 124166
rect 202420 124102 202472 124108
rect 202432 123622 202460 124102
rect 202420 123616 202472 123622
rect 202420 123558 202472 123564
rect 202328 123548 202380 123554
rect 202328 123490 202380 123496
rect 202340 114481 202368 123490
rect 202432 115841 202460 123558
rect 202892 122834 202920 124510
rect 203156 124432 203208 124438
rect 203156 124374 203208 124380
rect 203064 124296 203116 124302
rect 203064 124238 203116 124244
rect 202708 122806 202920 122834
rect 202972 122868 203024 122874
rect 202972 122810 203024 122816
rect 202708 122754 202736 122806
rect 202708 122726 202920 122754
rect 202892 117978 202920 122726
rect 202880 117972 202932 117978
rect 202880 117914 202932 117920
rect 202984 116618 203012 122810
rect 202972 116612 203024 116618
rect 202972 116554 203024 116560
rect 202418 115832 202474 115841
rect 202418 115767 202474 115776
rect 202326 114472 202382 114481
rect 202326 114407 202382 114416
rect 202236 113144 202288 113150
rect 202236 113086 202288 113092
rect 202050 111208 202106 111217
rect 202050 111143 202106 111152
rect 201866 109848 201922 109857
rect 201866 109783 201868 109792
rect 201920 109783 201922 109792
rect 201868 109754 201920 109760
rect 202248 106457 202276 113086
rect 202788 110424 202840 110430
rect 202788 110366 202840 110372
rect 202800 109177 202828 110366
rect 202786 109168 202842 109177
rect 202786 109103 202842 109112
rect 202788 107636 202840 107642
rect 202788 107578 202840 107584
rect 202800 107137 202828 107578
rect 202786 107128 202842 107137
rect 202786 107063 202842 107072
rect 202234 106448 202290 106457
rect 202234 106383 202290 106392
rect 201868 105596 201920 105602
rect 201868 105538 201920 105544
rect 201774 105088 201830 105097
rect 201774 105023 201830 105032
rect 201880 103737 201908 105538
rect 201866 103728 201922 103737
rect 201866 103663 201922 103672
rect 201880 103514 201908 103663
rect 201788 103486 201908 103514
rect 201682 103048 201738 103057
rect 201682 102983 201738 102992
rect 201590 100328 201646 100337
rect 201590 100263 201646 100272
rect 201604 100026 201632 100263
rect 201592 100020 201644 100026
rect 201592 99962 201644 99968
rect 201592 99340 201644 99346
rect 201592 99282 201644 99288
rect 201604 98977 201632 99282
rect 201590 98968 201646 98977
rect 201590 98903 201646 98912
rect 201788 98818 201816 103486
rect 201866 101688 201922 101697
rect 201866 101623 201922 101632
rect 201604 98790 201816 98818
rect 201498 82920 201554 82929
rect 201498 82855 201554 82864
rect 200670 77344 200726 77353
rect 200670 77279 200726 77288
rect 200486 75168 200542 75177
rect 200486 75103 200542 75112
rect 200500 74594 200528 75103
rect 200488 74588 200540 74594
rect 200488 74530 200540 74536
rect 200396 71664 200448 71670
rect 200396 71606 200448 71612
rect 200500 71482 200528 74530
rect 200578 73264 200634 73273
rect 200578 73199 200634 73208
rect 200408 71454 200528 71482
rect 200408 70174 200436 71454
rect 200488 71392 200540 71398
rect 200488 71334 200540 71340
rect 200396 70168 200448 70174
rect 200396 70110 200448 70116
rect 200500 70038 200528 71334
rect 200488 70032 200540 70038
rect 200488 69974 200540 69980
rect 200210 67416 200266 67425
rect 200592 67386 200620 73199
rect 200684 67590 200712 77279
rect 201314 76528 201370 76537
rect 201314 76463 201370 76472
rect 201328 75954 201356 76463
rect 201316 75948 201368 75954
rect 201316 75890 201368 75896
rect 200948 75880 201000 75886
rect 200948 75822 201000 75828
rect 200960 74769 200988 75822
rect 200946 74760 201002 74769
rect 200946 74695 201002 74704
rect 200854 73808 200910 73817
rect 200854 73743 200910 73752
rect 200762 72448 200818 72457
rect 200762 72383 200818 72392
rect 200672 67584 200724 67590
rect 200672 67526 200724 67532
rect 200210 67351 200266 67360
rect 200580 67380 200632 67386
rect 200580 67322 200632 67328
rect 199660 66972 199712 66978
rect 199660 66914 199712 66920
rect 198740 66904 198792 66910
rect 198740 66846 198792 66852
rect 200776 66026 200804 72383
rect 200868 66201 200896 73743
rect 201328 71398 201356 75890
rect 201512 71602 201540 82855
rect 201500 71596 201552 71602
rect 201500 71538 201552 71544
rect 201316 71392 201368 71398
rect 201316 71334 201368 71340
rect 201604 69766 201632 98790
rect 201880 98546 201908 101623
rect 202788 100088 202840 100094
rect 202788 100030 202840 100036
rect 202800 99657 202828 100030
rect 202786 99648 202842 99657
rect 202786 99583 202842 99592
rect 201696 98518 201908 98546
rect 201696 69902 201724 98518
rect 201958 97608 202014 97617
rect 201958 97543 202014 97552
rect 201776 90840 201828 90846
rect 201774 90808 201776 90817
rect 201828 90808 201830 90817
rect 201774 90743 201830 90752
rect 201774 90128 201830 90137
rect 201774 90063 201776 90072
rect 201828 90063 201830 90072
rect 201776 90034 201828 90040
rect 201972 89714 202000 97543
rect 202142 96520 202198 96529
rect 202142 96455 202198 96464
rect 202156 95946 202184 96455
rect 202418 96248 202474 96257
rect 202418 96183 202474 96192
rect 202144 95940 202196 95946
rect 202144 95882 202196 95888
rect 202050 92168 202106 92177
rect 202050 92103 202106 92112
rect 201788 89686 202000 89714
rect 201788 69970 201816 89686
rect 202064 84946 202092 92103
rect 202142 89448 202198 89457
rect 202142 89383 202198 89392
rect 201880 84918 202092 84946
rect 201880 71534 201908 84918
rect 202050 80608 202106 80617
rect 202050 80543 202106 80552
rect 201960 74520 202012 74526
rect 201960 74462 202012 74468
rect 201972 73817 202000 74462
rect 201958 73808 202014 73817
rect 201958 73743 202014 73752
rect 201960 71732 202012 71738
rect 201960 71674 202012 71680
rect 201868 71528 201920 71534
rect 201868 71470 201920 71476
rect 201972 71233 202000 71674
rect 201958 71224 202014 71233
rect 201958 71159 202014 71168
rect 202064 70553 202092 80543
rect 202050 70544 202106 70553
rect 202050 70479 202106 70488
rect 201776 69964 201828 69970
rect 201776 69906 201828 69912
rect 201684 69896 201736 69902
rect 201684 69838 201736 69844
rect 201592 69760 201644 69766
rect 201592 69702 201644 69708
rect 202156 69698 202184 89383
rect 202234 81968 202290 81977
rect 202234 81903 202290 81912
rect 202248 69834 202276 81903
rect 202236 69828 202288 69834
rect 202236 69770 202288 69776
rect 202144 69692 202196 69698
rect 202144 69634 202196 69640
rect 202432 69562 202460 96183
rect 203076 95946 203104 124238
rect 203168 109818 203196 124374
rect 203248 122936 203300 122942
rect 203248 122878 203300 122884
rect 203260 115258 203288 122878
rect 203248 115252 203300 115258
rect 203248 115194 203300 115200
rect 203156 109812 203208 109818
rect 203156 109754 203208 109760
rect 203064 95940 203116 95946
rect 203064 95882 203116 95888
rect 202788 94512 202840 94518
rect 202788 94454 202840 94460
rect 202800 94217 202828 94454
rect 202786 94208 202842 94217
rect 202786 94143 202842 94152
rect 202512 89684 202564 89690
rect 202512 89626 202564 89632
rect 202524 88777 202552 89626
rect 202510 88768 202566 88777
rect 202510 88703 202566 88712
rect 202512 88324 202564 88330
rect 202512 88266 202564 88272
rect 202524 88097 202552 88266
rect 202510 88088 202566 88097
rect 202510 88023 202566 88032
rect 202512 86964 202564 86970
rect 202512 86906 202564 86912
rect 202524 86737 202552 86906
rect 202510 86728 202566 86737
rect 202510 86663 202566 86672
rect 202696 84856 202748 84862
rect 202694 84824 202696 84833
rect 203248 84856 203300 84862
rect 202748 84824 202750 84833
rect 203248 84798 203300 84804
rect 202694 84759 202750 84768
rect 202694 84280 202750 84289
rect 202694 84215 202696 84224
rect 202748 84215 202750 84224
rect 203064 84244 203116 84250
rect 202696 84186 202748 84192
rect 203064 84186 203116 84192
rect 202510 80200 202566 80209
rect 202510 80135 202566 80144
rect 202524 69737 202552 80135
rect 202788 79348 202840 79354
rect 202788 79290 202840 79296
rect 202800 79257 202828 79290
rect 202786 79248 202842 79257
rect 202786 79183 202842 79192
rect 202788 78736 202840 78742
rect 202786 78704 202788 78713
rect 202840 78704 202842 78713
rect 202786 78639 202842 78648
rect 202510 69728 202566 69737
rect 202510 69663 202566 69672
rect 202788 69692 202840 69698
rect 202788 69634 202840 69640
rect 202420 69556 202472 69562
rect 202420 69498 202472 69504
rect 202696 69488 202748 69494
rect 202696 69430 202748 69436
rect 202604 68944 202656 68950
rect 202604 68886 202656 68892
rect 202616 68338 202644 68886
rect 202708 68678 202736 69430
rect 202800 69018 202828 69634
rect 202788 69012 202840 69018
rect 202788 68954 202840 68960
rect 202696 68672 202748 68678
rect 202696 68614 202748 68620
rect 202604 68332 202656 68338
rect 202604 68274 202656 68280
rect 200854 66192 200910 66201
rect 200854 66127 200910 66136
rect 200764 66020 200816 66026
rect 200764 65962 200816 65968
rect 203076 65550 203104 84186
rect 203156 83496 203208 83502
rect 203156 83438 203208 83444
rect 203168 83337 203196 83438
rect 203154 83328 203210 83337
rect 203154 83263 203210 83272
rect 203168 65958 203196 83263
rect 203260 70242 203288 84798
rect 203340 79348 203392 79354
rect 203340 79290 203392 79296
rect 203248 70236 203300 70242
rect 203248 70178 203300 70184
rect 203156 65952 203208 65958
rect 203156 65894 203208 65900
rect 203352 65618 203380 79290
rect 203444 67182 203472 168302
rect 203708 121916 203760 121922
rect 203708 121858 203760 121864
rect 203616 120556 203668 120562
rect 203616 120498 203668 120504
rect 203524 120488 203576 120494
rect 203524 120430 203576 120436
rect 203432 67176 203484 67182
rect 203432 67118 203484 67124
rect 203340 65612 203392 65618
rect 203340 65554 203392 65560
rect 203064 65544 203116 65550
rect 203064 65486 203116 65492
rect 198648 21412 198700 21418
rect 198648 21354 198700 21360
rect 188344 18624 188396 18630
rect 188344 18566 188396 18572
rect 187608 5024 187660 5030
rect 187608 4966 187660 4972
rect 203536 3602 203564 120430
rect 203628 60722 203656 120498
rect 203720 102814 203748 121858
rect 203708 102808 203760 102814
rect 203708 102750 203760 102756
rect 204180 68338 204208 169934
rect 204352 167612 204404 167618
rect 204352 167554 204404 167560
rect 204364 69850 204392 167554
rect 204628 123208 204680 123214
rect 204628 123150 204680 123156
rect 204536 123072 204588 123078
rect 204536 123014 204588 123020
rect 204442 122904 204498 122913
rect 204442 122839 204498 122848
rect 204456 90846 204484 122839
rect 204548 94518 204576 123014
rect 204640 100026 204668 123150
rect 204720 123004 204772 123010
rect 204720 122946 204772 122952
rect 204732 110430 204760 122946
rect 204720 110424 204772 110430
rect 204720 110366 204772 110372
rect 204732 109750 204760 110366
rect 204720 109744 204772 109750
rect 204720 109686 204772 109692
rect 204628 100020 204680 100026
rect 204628 99962 204680 99968
rect 204536 94512 204588 94518
rect 204536 94454 204588 94460
rect 204444 90840 204496 90846
rect 204444 90782 204496 90788
rect 204456 90370 204484 90782
rect 204444 90364 204496 90370
rect 204444 90306 204496 90312
rect 204444 78736 204496 78742
rect 204444 78678 204496 78684
rect 204456 70310 204484 78678
rect 204824 70718 204852 169934
rect 205732 123412 205784 123418
rect 205732 123354 205784 123360
rect 205744 107642 205772 123354
rect 205732 107636 205784 107642
rect 205732 107578 205784 107584
rect 204812 70712 204864 70718
rect 204812 70654 204864 70660
rect 204444 70304 204496 70310
rect 204444 70246 204496 70252
rect 204364 69822 204484 69850
rect 204168 68332 204220 68338
rect 204168 68274 204220 68280
rect 204456 67590 204484 69822
rect 206112 69494 206140 169934
rect 207400 169318 207428 169934
rect 207388 169312 207440 169318
rect 207388 169254 207440 169260
rect 208688 169046 208716 169934
rect 208676 169040 208728 169046
rect 208676 168982 208728 168988
rect 209688 169040 209740 169046
rect 209688 168982 209740 168988
rect 209700 167346 209728 168982
rect 209688 167340 209740 167346
rect 209688 167282 209740 167288
rect 209044 165028 209096 165034
rect 209044 164970 209096 164976
rect 209056 124166 209084 164970
rect 208400 124160 208452 124166
rect 208400 124102 208452 124108
rect 209044 124160 209096 124166
rect 209044 124102 209096 124108
rect 208412 123350 208440 124102
rect 208400 123344 208452 123350
rect 208400 123286 208452 123292
rect 206284 121780 206336 121786
rect 206284 121722 206336 121728
rect 206100 69488 206152 69494
rect 206100 69430 206152 69436
rect 204444 67584 204496 67590
rect 204444 67526 204496 67532
rect 204456 67318 204484 67526
rect 204444 67312 204496 67318
rect 204444 67254 204496 67260
rect 203616 60716 203668 60722
rect 203616 60658 203668 60664
rect 206296 7614 206324 121722
rect 208412 100094 208440 123286
rect 208400 100088 208452 100094
rect 208400 100030 208452 100036
rect 208400 90092 208452 90098
rect 208400 90034 208452 90040
rect 208412 66230 208440 90034
rect 210620 69698 210648 169934
rect 211908 71058 211936 169934
rect 211896 71052 211948 71058
rect 211896 70994 211948 71000
rect 210608 69692 210660 69698
rect 210608 69634 210660 69640
rect 212552 69018 212580 169934
rect 213840 169386 213868 169934
rect 215128 169522 215156 169934
rect 215116 169516 215168 169522
rect 215116 169458 215168 169464
rect 213828 169380 213880 169386
rect 213828 169322 213880 169328
rect 215208 166388 215260 166394
rect 215208 166330 215260 166336
rect 215220 84862 215248 166330
rect 215208 84856 215260 84862
rect 215208 84798 215260 84804
rect 212540 69012 212592 69018
rect 212540 68954 212592 68960
rect 213828 69012 213880 69018
rect 213828 68954 213880 68960
rect 213840 68406 213868 68954
rect 213828 68400 213880 68406
rect 213828 68342 213880 68348
rect 215300 67516 215352 67522
rect 215300 67458 215352 67464
rect 215312 66910 215340 67458
rect 216416 66910 216444 169934
rect 217060 168026 217088 169934
rect 218348 168201 218376 169934
rect 218334 168192 218390 168201
rect 218334 168127 218336 168136
rect 218388 168127 218390 168136
rect 218336 168098 218388 168104
rect 218348 168067 218376 168098
rect 219636 168094 219664 169934
rect 220280 168230 220308 169934
rect 221568 169697 221596 169934
rect 221554 169688 221610 169697
rect 221554 169623 221610 169632
rect 221568 168230 221596 169623
rect 220268 168224 220320 168230
rect 220268 168166 220320 168172
rect 221556 168224 221608 168230
rect 221556 168166 221608 168172
rect 219624 168088 219676 168094
rect 219624 168030 219676 168036
rect 217048 168020 217100 168026
rect 217048 167962 217100 167968
rect 221568 166994 221596 168166
rect 221476 166966 221596 166994
rect 217968 159384 218020 159390
rect 217968 159326 218020 159332
rect 217980 79354 218008 159326
rect 220728 131776 220780 131782
rect 220728 131718 220780 131724
rect 220740 129062 220768 131718
rect 219440 129056 219492 129062
rect 219440 128998 219492 129004
rect 220728 129056 220780 129062
rect 220728 128998 220780 129004
rect 219452 99346 219480 128998
rect 220084 121712 220136 121718
rect 220084 121654 220136 121660
rect 219440 99340 219492 99346
rect 219440 99282 219492 99288
rect 217968 79348 218020 79354
rect 217968 79290 218020 79296
rect 215300 66904 215352 66910
rect 215300 66846 215352 66852
rect 216404 66904 216456 66910
rect 216404 66846 216456 66852
rect 208400 66224 208452 66230
rect 208400 66166 208452 66172
rect 208412 65754 208440 66166
rect 208400 65748 208452 65754
rect 208400 65690 208452 65696
rect 209044 65748 209096 65754
rect 209044 65690 209096 65696
rect 209056 17270 209084 65690
rect 220096 22778 220124 121654
rect 221476 74526 221504 166966
rect 222856 75886 222884 169934
rect 224788 167550 224816 169934
rect 226076 168366 226104 169934
rect 226064 168360 226116 168366
rect 226064 168302 226116 168308
rect 226076 167793 226104 168302
rect 227364 167958 227392 169934
rect 228744 168298 228772 170326
rect 228732 168292 228784 168298
rect 228732 168234 228784 168240
rect 227352 167952 227404 167958
rect 227352 167894 227404 167900
rect 226062 167784 226118 167793
rect 226062 167719 226118 167728
rect 224776 167544 224828 167550
rect 224776 167486 224828 167492
rect 226984 166456 227036 166462
rect 226984 166398 227036 166404
rect 224868 163600 224920 163606
rect 224868 163542 224920 163548
rect 224880 83502 224908 163542
rect 226340 122120 226392 122126
rect 226340 122062 226392 122068
rect 226352 121718 226380 122062
rect 226996 121718 227024 166398
rect 228836 161474 228864 170342
rect 228744 161446 228864 161474
rect 229112 170326 229310 170354
rect 226340 121712 226392 121718
rect 226340 121654 226392 121660
rect 226984 121712 227036 121718
rect 226984 121654 227036 121660
rect 226352 88330 226380 121654
rect 227720 120896 227772 120902
rect 227720 120838 227772 120844
rect 227732 120426 227760 120838
rect 228744 120426 228772 161446
rect 229112 159390 229140 170326
rect 229282 169552 229338 169561
rect 229282 169487 229338 169496
rect 229296 169114 229324 169487
rect 229284 169108 229336 169114
rect 229284 169050 229336 169056
rect 229388 165374 229416 196143
rect 229466 195392 229522 195401
rect 229466 195327 229522 195336
rect 229376 165368 229428 165374
rect 229376 165310 229428 165316
rect 229480 164898 229508 195327
rect 229558 192808 229614 192817
rect 229558 192743 229614 192752
rect 229572 165442 229600 192743
rect 229560 165436 229612 165442
rect 229560 165378 229612 165384
rect 229468 164892 229520 164898
rect 229468 164834 229520 164840
rect 229100 159384 229152 159390
rect 229100 159326 229152 159332
rect 229664 123690 229692 226306
rect 229848 209774 229876 228919
rect 230032 219065 230060 241538
rect 230124 221105 230152 242966
rect 230216 225865 230244 245618
rect 230308 227225 230336 247046
rect 230940 244452 230992 244458
rect 230940 244394 230992 244400
rect 230756 237516 230808 237522
rect 230756 237458 230808 237464
rect 230572 236020 230624 236026
rect 230572 235962 230624 235968
rect 230480 234660 230532 234666
rect 230480 234602 230532 234608
rect 230388 233300 230440 233306
rect 230388 233242 230440 233248
rect 230294 227216 230350 227225
rect 230294 227151 230350 227160
rect 230202 225856 230258 225865
rect 230202 225791 230258 225800
rect 230110 221096 230166 221105
rect 230110 221031 230166 221040
rect 230018 219056 230074 219065
rect 230018 218991 230074 219000
rect 230400 209778 230428 233242
rect 230492 210905 230520 234602
rect 230584 212945 230612 235962
rect 230664 230852 230716 230858
rect 230664 230794 230716 230800
rect 230570 212936 230626 212945
rect 230570 212871 230626 212880
rect 230570 212256 230626 212265
rect 230570 212191 230626 212200
rect 230478 210896 230534 210905
rect 230478 210831 230534 210840
rect 229848 209746 229968 209774
rect 229836 208412 229888 208418
rect 229836 208354 229888 208360
rect 229848 200114 229876 208354
rect 229940 204105 229968 209746
rect 230388 209772 230440 209778
rect 230388 209714 230440 209720
rect 230400 209545 230428 209714
rect 230386 209536 230442 209545
rect 230386 209471 230442 209480
rect 230400 208418 230428 209471
rect 230388 208412 230440 208418
rect 230388 208354 230440 208360
rect 230018 207496 230074 207505
rect 230018 207431 230074 207440
rect 229926 204096 229982 204105
rect 229926 204031 229982 204040
rect 229848 200086 229968 200114
rect 229742 181112 229798 181121
rect 229742 181047 229798 181056
rect 229652 123684 229704 123690
rect 229652 123626 229704 123632
rect 229756 123486 229784 181047
rect 229100 123480 229152 123486
rect 229100 123422 229152 123428
rect 229744 123480 229796 123486
rect 229744 123422 229796 123428
rect 227720 120420 227772 120426
rect 227720 120362 227772 120368
rect 228732 120420 228784 120426
rect 228732 120362 228784 120368
rect 227732 93854 227760 120362
rect 227732 93826 227852 93854
rect 226340 88324 226392 88330
rect 226340 88266 226392 88272
rect 226800 88324 226852 88330
rect 226800 88266 226852 88272
rect 226812 87650 226840 88266
rect 226800 87644 226852 87650
rect 226800 87586 226852 87592
rect 227824 86970 227852 93826
rect 229112 89690 229140 123422
rect 229940 113150 229968 200086
rect 230032 166326 230060 207431
rect 230020 166320 230072 166326
rect 230020 166262 230072 166268
rect 229928 113144 229980 113150
rect 229928 113086 229980 113092
rect 230492 107642 230520 210831
rect 230584 109002 230612 212191
rect 230676 206145 230704 230794
rect 230768 214305 230796 237458
rect 230848 229152 230900 229158
rect 230848 229094 230900 229100
rect 230754 214296 230810 214305
rect 230754 214231 230810 214240
rect 230662 206136 230718 206145
rect 230662 206071 230718 206080
rect 230572 108996 230624 109002
rect 230572 108938 230624 108944
rect 230480 107636 230532 107642
rect 230480 107578 230532 107584
rect 230676 105602 230704 206071
rect 230860 160750 230888 229094
rect 230952 223582 230980 244394
rect 231308 244384 231360 244390
rect 231308 244326 231360 244332
rect 231032 241528 231084 241534
rect 231032 241470 231084 241476
rect 231044 229090 231072 241470
rect 231216 238808 231268 238814
rect 231216 238750 231268 238756
rect 231124 237448 231176 237454
rect 231124 237390 231176 237396
rect 231032 229084 231084 229090
rect 231032 229026 231084 229032
rect 230940 223576 230992 223582
rect 230940 223518 230992 223524
rect 230952 222465 230980 223518
rect 230938 222456 230994 222465
rect 230938 222391 230994 222400
rect 230952 164966 230980 222391
rect 231136 215665 231164 237390
rect 231228 217025 231256 238750
rect 231320 223825 231348 244326
rect 231952 242956 232004 242962
rect 231952 242898 232004 242904
rect 231964 230450 231992 242898
rect 232688 236768 232740 236774
rect 232688 236710 232740 236716
rect 231952 230444 232004 230450
rect 231952 230386 232004 230392
rect 232320 229900 232372 229906
rect 232320 229842 232372 229848
rect 231952 229764 232004 229770
rect 231952 229706 232004 229712
rect 231860 229220 231912 229226
rect 231860 229162 231912 229168
rect 231400 229084 231452 229090
rect 231400 229026 231452 229032
rect 231306 223816 231362 223825
rect 231306 223751 231362 223760
rect 231412 220425 231440 229026
rect 231398 220416 231454 220425
rect 231398 220351 231454 220360
rect 231412 219434 231440 220351
rect 231320 219406 231440 219434
rect 231214 217016 231270 217025
rect 231214 216951 231270 216960
rect 231122 215656 231178 215665
rect 231122 215591 231178 215600
rect 231030 174856 231086 174865
rect 231030 174791 231086 174800
rect 230940 164960 230992 164966
rect 230940 164902 230992 164908
rect 231044 163538 231072 174791
rect 231032 163532 231084 163538
rect 231032 163474 231084 163480
rect 230848 160744 230900 160750
rect 230848 160686 230900 160692
rect 231320 142866 231348 219406
rect 231872 185065 231900 229162
rect 231858 185056 231914 185065
rect 231858 184991 231914 185000
rect 231858 179616 231914 179625
rect 231858 179551 231914 179560
rect 231766 171864 231822 171873
rect 231766 171799 231768 171808
rect 231820 171799 231822 171808
rect 231768 171770 231820 171776
rect 231674 171184 231730 171193
rect 231674 171119 231730 171128
rect 231688 171086 231716 171119
rect 231676 171080 231728 171086
rect 231676 171022 231728 171028
rect 231780 170218 231808 171770
rect 231872 170406 231900 179551
rect 231964 176225 231992 229706
rect 232136 229696 232188 229702
rect 232136 229638 232188 229644
rect 232044 229356 232096 229362
rect 232044 229298 232096 229304
rect 232056 178265 232084 229298
rect 232148 184385 232176 229638
rect 232228 229628 232280 229634
rect 232228 229570 232280 229576
rect 232240 189825 232268 229570
rect 232332 192545 232360 229842
rect 232504 229560 232556 229566
rect 232504 229502 232556 229508
rect 232412 229492 232464 229498
rect 232412 229434 232464 229440
rect 232424 194585 232452 229434
rect 232516 200114 232544 229502
rect 232596 229424 232648 229430
rect 232596 229366 232648 229372
rect 232608 200705 232636 229366
rect 232700 225185 232728 236710
rect 233240 232008 233292 232014
rect 233240 231950 233292 231956
rect 232686 225176 232742 225185
rect 232686 225111 232742 225120
rect 232688 218000 232740 218006
rect 232686 217968 232688 217977
rect 232740 217968 232742 217977
rect 232686 217903 232742 217912
rect 232686 206136 232742 206145
rect 232686 206071 232742 206080
rect 232700 205698 232728 206071
rect 232688 205692 232740 205698
rect 232688 205634 232740 205640
rect 233146 204776 233202 204785
rect 233146 204711 233202 204720
rect 233160 204338 233188 204711
rect 233148 204332 233200 204338
rect 233148 204274 233200 204280
rect 232688 204264 232740 204270
rect 232688 204206 232740 204212
rect 232700 204105 232728 204206
rect 232686 204096 232742 204105
rect 232686 204031 232742 204040
rect 232688 202836 232740 202842
rect 232688 202778 232740 202784
rect 232700 202745 232728 202778
rect 232686 202736 232742 202745
rect 232686 202671 232742 202680
rect 232594 200696 232650 200705
rect 232594 200631 232650 200640
rect 232516 200086 232728 200114
rect 232700 199345 232728 200086
rect 232686 199336 232742 199345
rect 232686 199271 232742 199280
rect 232594 197976 232650 197985
rect 232594 197911 232650 197920
rect 232410 194576 232466 194585
rect 232410 194511 232466 194520
rect 232318 192536 232374 192545
rect 232318 192471 232374 192480
rect 232226 189816 232282 189825
rect 232226 189751 232282 189760
rect 232134 184376 232190 184385
rect 232134 184311 232190 184320
rect 232410 183016 232466 183025
rect 232410 182951 232466 182960
rect 232226 180296 232282 180305
rect 232226 180231 232282 180240
rect 232042 178256 232098 178265
rect 232042 178191 232098 178200
rect 231950 176216 232006 176225
rect 231950 176151 232006 176160
rect 232042 173496 232098 173505
rect 232042 173431 232098 173440
rect 231952 171080 232004 171086
rect 231952 171022 232004 171028
rect 231860 170400 231912 170406
rect 231860 170342 231912 170348
rect 231780 170190 231900 170218
rect 231872 165306 231900 170190
rect 231860 165300 231912 165306
rect 231860 165242 231912 165248
rect 231964 165102 231992 171022
rect 231952 165096 232004 165102
rect 231952 165038 232004 165044
rect 232056 163606 232084 173431
rect 232240 166462 232268 180231
rect 232228 166456 232280 166462
rect 232228 166398 232280 166404
rect 232424 165510 232452 182951
rect 232502 176896 232558 176905
rect 232502 176831 232558 176840
rect 232516 166394 232544 176831
rect 232504 166388 232556 166394
rect 232504 166330 232556 166336
rect 232412 165504 232464 165510
rect 232412 165446 232464 165452
rect 232044 163600 232096 163606
rect 232044 163542 232096 163548
rect 231308 142860 231360 142866
rect 231308 142802 231360 142808
rect 232608 131782 232636 197911
rect 232700 165034 232728 199271
rect 233146 191176 233202 191185
rect 233146 191111 233148 191120
rect 233200 191111 233202 191120
rect 233148 191082 233200 191088
rect 232778 188456 232834 188465
rect 232778 188391 232834 188400
rect 232792 165170 232820 188391
rect 233148 188352 233200 188358
rect 233148 188294 233200 188300
rect 233160 187785 233188 188294
rect 233146 187776 233202 187785
rect 233146 187711 233202 187720
rect 233148 186992 233200 186998
rect 233148 186934 233200 186940
rect 233160 186425 233188 186934
rect 233146 186416 233202 186425
rect 233146 186351 233202 186360
rect 233056 175228 233108 175234
rect 233056 175170 233108 175176
rect 233068 174865 233096 175170
rect 233054 174856 233110 174865
rect 233054 174791 233110 174800
rect 233252 167754 233280 231950
rect 233896 218006 233924 683130
rect 233976 563100 234028 563106
rect 233976 563042 234028 563048
rect 233988 229090 234016 563042
rect 234068 351960 234120 351966
rect 234068 351902 234120 351908
rect 233976 229084 234028 229090
rect 233976 229026 234028 229032
rect 233884 218000 233936 218006
rect 233884 217942 233936 217948
rect 234080 209778 234108 351902
rect 234632 256018 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 700534 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 267648 700528 267700 700534
rect 267648 700470 267700 700476
rect 249064 643136 249116 643142
rect 249064 643078 249116 643084
rect 239404 630692 239456 630698
rect 239404 630634 239456 630640
rect 235264 616888 235316 616894
rect 235264 616830 235316 616836
rect 234620 256012 234672 256018
rect 234620 255954 234672 255960
rect 234620 232076 234672 232082
rect 234620 232018 234672 232024
rect 234068 209772 234120 209778
rect 234068 209714 234120 209720
rect 233330 201376 233386 201385
rect 233330 201311 233386 201320
rect 233344 200802 233372 201311
rect 233332 200796 233384 200802
rect 233332 200738 233384 200744
rect 233240 167748 233292 167754
rect 233240 167690 233292 167696
rect 233344 166977 233372 200738
rect 233884 191888 233936 191894
rect 233884 191830 233936 191836
rect 233424 191140 233476 191146
rect 233424 191082 233476 191088
rect 233330 166968 233386 166977
rect 233330 166903 233386 166912
rect 233436 165578 233464 191082
rect 233516 188352 233568 188358
rect 233516 188294 233568 188300
rect 233424 165572 233476 165578
rect 233424 165514 233476 165520
rect 233528 165238 233556 188294
rect 233608 186992 233660 186998
rect 233608 186934 233660 186940
rect 233620 165617 233648 186934
rect 233896 170105 233924 191830
rect 233882 170096 233938 170105
rect 233882 170031 233938 170040
rect 233606 165608 233662 165617
rect 233606 165543 233662 165552
rect 233516 165232 233568 165238
rect 233516 165174 233568 165180
rect 232780 165164 232832 165170
rect 232780 165106 232832 165112
rect 232688 165028 232740 165034
rect 232688 164970 232740 164976
rect 232596 131776 232648 131782
rect 232596 131718 232648 131724
rect 234632 126954 234660 232018
rect 234712 231872 234764 231878
rect 234712 231814 234764 231820
rect 234724 167686 234752 231814
rect 235276 169454 235304 616830
rect 238024 378208 238076 378214
rect 238024 378150 238076 378156
rect 235356 230648 235408 230654
rect 235356 230590 235408 230596
rect 235368 219434 235396 230590
rect 235356 219428 235408 219434
rect 235356 219370 235408 219376
rect 238036 169590 238064 378150
rect 238024 169584 238076 169590
rect 238024 169526 238076 169532
rect 235264 169448 235316 169454
rect 235264 169390 235316 169396
rect 239416 168162 239444 630634
rect 242164 590708 242216 590714
rect 242164 590650 242216 590656
rect 242176 188358 242204 590650
rect 244924 364404 244976 364410
rect 244924 364346 244976 364352
rect 242164 188352 242216 188358
rect 242164 188294 242216 188300
rect 239404 168156 239456 168162
rect 239404 168098 239456 168104
rect 234712 167680 234764 167686
rect 234712 167622 234764 167628
rect 244936 167482 244964 364346
rect 249076 186998 249104 643078
rect 278044 536852 278096 536858
rect 278044 536794 278096 536800
rect 278056 204270 278084 536794
rect 282932 239426 282960 702406
rect 289084 470620 289136 470626
rect 289084 470562 289136 470568
rect 282920 239420 282972 239426
rect 282920 239362 282972 239368
rect 278044 204264 278096 204270
rect 278044 204206 278096 204212
rect 289096 202842 289124 470562
rect 289084 202836 289136 202842
rect 289084 202778 289136 202784
rect 249064 186992 249116 186998
rect 249064 186934 249116 186940
rect 299492 168230 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 331232 233238 331260 702986
rect 348804 702434 348832 703520
rect 347792 702406 348832 702434
rect 331220 233232 331272 233238
rect 331220 233174 331272 233180
rect 347792 168366 347820 702406
rect 364996 700466 365024 703520
rect 364984 700460 365036 700466
rect 364984 700402 365036 700408
rect 397472 699718 397500 703520
rect 396724 699712 396776 699718
rect 396724 699654 396776 699660
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 396736 168910 396764 699654
rect 412652 232558 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 429856 700398 429884 703520
rect 429844 700392 429896 700398
rect 429844 700334 429896 700340
rect 412640 232552 412692 232558
rect 412640 232494 412692 232500
rect 462332 171834 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 477512 200802 477540 702406
rect 477500 200796 477552 200802
rect 477500 200738 477552 200744
rect 494072 175234 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 700330 527220 703520
rect 543476 702434 543504 703520
rect 559668 702434 559696 703520
rect 542372 702406 543504 702434
rect 558932 702406 559696 702434
rect 527180 700324 527232 700330
rect 527180 700266 527232 700272
rect 542372 257378 542400 702406
rect 542360 257372 542412 257378
rect 542360 257314 542412 257320
rect 548616 226364 548668 226370
rect 548616 226306 548668 226312
rect 548628 206990 548656 226306
rect 558932 223582 558960 702406
rect 580262 697232 580318 697241
rect 580262 697167 580318 697176
rect 579618 683904 579674 683913
rect 579618 683839 579674 683848
rect 579632 683194 579660 683839
rect 579620 683188 579672 683194
rect 579620 683130 579672 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 579894 537840 579950 537849
rect 579894 537775 579950 537784
rect 579908 536858 579936 537775
rect 579896 536852 579948 536858
rect 579896 536794 579948 536800
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580184 470626 580212 471407
rect 580172 470620 580224 470626
rect 580172 470562 580224 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 579802 365120 579858 365129
rect 579802 365055 579858 365064
rect 579816 364410 579844 365055
rect 579804 364404 579856 364410
rect 579804 364346 579856 364352
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 579618 325272 579674 325281
rect 579618 325207 579674 325216
rect 579632 324358 579660 325207
rect 579620 324352 579672 324358
rect 579620 324294 579672 324300
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 311914 580212 312015
rect 580172 311908 580224 311914
rect 580172 311850 580224 311856
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 578882 272232 578938 272241
rect 578882 272167 578938 272176
rect 558920 223576 558972 223582
rect 558920 223518 558972 223524
rect 548616 206984 548668 206990
rect 548616 206926 548668 206932
rect 548524 205692 548576 205698
rect 548524 205634 548576 205640
rect 494060 175228 494112 175234
rect 494060 175170 494112 175176
rect 462320 171828 462372 171834
rect 462320 171770 462372 171776
rect 396724 168904 396776 168910
rect 396724 168846 396776 168852
rect 347780 168360 347832 168366
rect 347780 168302 347832 168308
rect 299480 168224 299532 168230
rect 299480 168166 299532 168172
rect 244924 167476 244976 167482
rect 244924 167418 244976 167424
rect 548536 167006 548564 205634
rect 578896 191146 578924 272167
rect 579986 258904 580042 258913
rect 579986 258839 580042 258848
rect 580000 258126 580028 258839
rect 579988 258120 580040 258126
rect 579988 258062 580040 258068
rect 580170 245576 580226 245585
rect 580170 245511 580226 245520
rect 580184 244322 580212 245511
rect 580172 244316 580224 244322
rect 580172 244258 580224 244264
rect 580276 233889 580304 697167
rect 580354 524512 580410 524521
rect 580354 524447 580410 524456
rect 580368 236706 580396 524447
rect 580446 431624 580502 431633
rect 580446 431559 580502 431568
rect 580356 236700 580408 236706
rect 580356 236642 580408 236648
rect 580262 233880 580318 233889
rect 580262 233815 580318 233824
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 580000 231130 580028 232319
rect 579988 231124 580040 231130
rect 579988 231066 580040 231072
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 579988 206984 580040 206990
rect 579988 206926 580040 206932
rect 580000 205737 580028 206926
rect 579986 205728 580042 205737
rect 579986 205663 580042 205672
rect 580264 204332 580316 204338
rect 580264 204274 580316 204280
rect 579710 192536 579766 192545
rect 579710 192471 579766 192480
rect 579724 191894 579752 192471
rect 579712 191888 579764 191894
rect 579712 191830 579764 191836
rect 578884 191140 578936 191146
rect 578884 191082 578936 191088
rect 580276 179217 580304 204274
rect 580262 179208 580318 179217
rect 580262 179143 580318 179152
rect 580460 169046 580488 431559
rect 580448 169040 580500 169046
rect 580448 168982 580500 168988
rect 548524 167000 548576 167006
rect 548524 166942 548576 166948
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580264 162172 580316 162178
rect 580264 162114 580316 162120
rect 580276 152697 580304 162114
rect 580262 152688 580318 152697
rect 580262 152623 580318 152632
rect 580262 139360 580318 139369
rect 580262 139295 580318 139304
rect 580276 127634 580304 139295
rect 580264 127628 580316 127634
rect 580264 127570 580316 127576
rect 234620 126948 234672 126954
rect 234620 126890 234672 126896
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 234632 126274 234660 126890
rect 234620 126268 234672 126274
rect 234620 126210 234672 126216
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 306380 124228 306432 124234
rect 306380 124170 306432 124176
rect 259460 123140 259512 123146
rect 259460 123082 259512 123088
rect 252560 120352 252612 120358
rect 252560 120294 252612 120300
rect 235264 120284 235316 120290
rect 235264 120226 235316 120232
rect 231768 108996 231820 109002
rect 231768 108938 231820 108944
rect 231780 108322 231808 108938
rect 231768 108316 231820 108322
rect 231768 108258 231820 108264
rect 231768 107636 231820 107642
rect 231768 107578 231820 107584
rect 231780 106962 231808 107578
rect 231768 106956 231820 106962
rect 231768 106898 231820 106904
rect 230664 105596 230716 105602
rect 230664 105538 230716 105544
rect 229100 89684 229152 89690
rect 229100 89626 229152 89632
rect 230388 89684 230440 89690
rect 230388 89626 230440 89632
rect 230400 89010 230428 89626
rect 230388 89004 230440 89010
rect 230388 88946 230440 88952
rect 227812 86964 227864 86970
rect 227812 86906 227864 86912
rect 227824 86290 227852 86906
rect 227812 86284 227864 86290
rect 227812 86226 227864 86232
rect 233884 85604 233936 85610
rect 233884 85546 233936 85552
rect 224868 83496 224920 83502
rect 224868 83438 224920 83444
rect 222844 75880 222896 75886
rect 222844 75822 222896 75828
rect 223488 75880 223540 75886
rect 223488 75822 223540 75828
rect 223500 75206 223528 75822
rect 223488 75200 223540 75206
rect 223488 75142 223540 75148
rect 221464 74520 221516 74526
rect 221464 74462 221516 74468
rect 233896 67590 233924 85546
rect 233884 67584 233936 67590
rect 233884 67526 233936 67532
rect 220084 22772 220136 22778
rect 220084 22714 220136 22720
rect 209044 17264 209096 17270
rect 209044 17206 209096 17212
rect 206284 7608 206336 7614
rect 206284 7550 206336 7556
rect 235276 3738 235304 120226
rect 251180 119468 251232 119474
rect 251180 119410 251232 119416
rect 238760 86284 238812 86290
rect 238760 86226 238812 86232
rect 238772 16574 238800 86226
rect 241520 79348 241572 79354
rect 241520 79290 241572 79296
rect 241532 16574 241560 79290
rect 249800 64388 249852 64394
rect 249800 64330 249852 64336
rect 242900 61532 242952 61538
rect 242900 61474 242952 61480
rect 238772 16546 239352 16574
rect 241532 16546 241744 16574
rect 235264 3732 235316 3738
rect 235264 3674 235316 3680
rect 203524 3596 203576 3602
rect 203524 3538 203576 3544
rect 184204 3528 184256 3534
rect 184204 3470 184256 3476
rect 177304 3460 177356 3466
rect 177304 3402 177356 3408
rect 239324 480 239352 16546
rect 240140 11756 240192 11762
rect 240140 11698 240192 11704
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240152 354 240180 11698
rect 241716 480 241744 16546
rect 242912 3670 242940 61474
rect 248420 60104 248472 60110
rect 248420 60046 248472 60052
rect 245660 49088 245712 49094
rect 245660 49030 245712 49036
rect 245672 16574 245700 49030
rect 247040 46232 247092 46238
rect 247040 46174 247092 46180
rect 247052 16574 247080 46174
rect 245672 16546 245976 16574
rect 247052 16546 247632 16574
rect 242992 7676 243044 7682
rect 242992 7618 243044 7624
rect 242900 3664 242952 3670
rect 242900 3606 242952 3612
rect 243004 3482 243032 7618
rect 245200 3800 245252 3806
rect 245200 3742 245252 3748
rect 244096 3664 244148 3670
rect 244096 3606 244148 3612
rect 242912 3454 243032 3482
rect 242912 480 242940 3454
rect 244108 480 244136 3606
rect 245212 480 245240 3742
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 247604 480 247632 16546
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248432 354 248460 60046
rect 249812 16574 249840 64330
rect 249812 16546 250024 16574
rect 249996 480 250024 16546
rect 251192 3670 251220 119410
rect 251272 50380 251324 50386
rect 251272 50322 251324 50328
rect 251180 3664 251232 3670
rect 251180 3606 251232 3612
rect 251284 3482 251312 50322
rect 252572 16574 252600 120294
rect 255320 102808 255372 102814
rect 255320 102750 255372 102756
rect 253940 75948 253992 75954
rect 253940 75890 253992 75896
rect 253952 16574 253980 75890
rect 255332 16574 255360 102750
rect 256700 100088 256752 100094
rect 256700 100030 256752 100036
rect 252572 16546 253520 16574
rect 253952 16546 254256 16574
rect 255332 16546 255912 16574
rect 252376 3664 252428 3670
rect 252376 3606 252428 3612
rect 251192 3454 251312 3482
rect 251192 480 251220 3454
rect 252388 480 252416 3606
rect 253492 480 253520 16546
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255884 480 255912 16546
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256712 354 256740 100030
rect 258724 99408 258776 99414
rect 258724 99350 258776 99356
rect 258736 67454 258764 99350
rect 258724 67448 258776 67454
rect 258724 67390 258776 67396
rect 258264 14476 258316 14482
rect 258264 14418 258316 14424
rect 258276 480 258304 14418
rect 259472 11762 259500 123082
rect 292580 122324 292632 122330
rect 292580 122266 292632 122272
rect 271880 119400 271932 119406
rect 271880 119342 271932 119348
rect 267832 109812 267884 109818
rect 267832 109754 267884 109760
rect 260840 95940 260892 95946
rect 260840 95882 260892 95888
rect 259552 61464 259604 61470
rect 259552 61406 259604 61412
rect 259460 11756 259512 11762
rect 259460 11698 259512 11704
rect 259564 6914 259592 61406
rect 260852 16574 260880 95882
rect 262220 62960 262272 62966
rect 262220 62902 262272 62908
rect 262232 16574 262260 62902
rect 264244 55956 264296 55962
rect 264244 55898 264296 55904
rect 263600 24132 263652 24138
rect 263600 24074 263652 24080
rect 263612 16574 263640 24074
rect 260852 16546 261800 16574
rect 262232 16546 262536 16574
rect 263612 16546 264192 16574
rect 260656 11756 260708 11762
rect 260656 11698 260708 11704
rect 259472 6886 259592 6914
rect 259472 480 259500 6886
rect 260668 480 260696 11698
rect 261772 480 261800 16546
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 264164 480 264192 16546
rect 264256 3194 264284 55898
rect 266360 21412 266412 21418
rect 266360 21354 266412 21360
rect 266372 16574 266400 21354
rect 267844 16574 267872 109754
rect 270500 64320 270552 64326
rect 270500 64262 270552 64268
rect 269120 39364 269172 39370
rect 269120 39306 269172 39312
rect 269132 16574 269160 39306
rect 270512 16574 270540 64262
rect 271892 16574 271920 119342
rect 282920 116612 282972 116618
rect 282920 116554 282972 116560
rect 277400 84856 277452 84862
rect 277400 84798 277452 84804
rect 273260 57248 273312 57254
rect 273260 57190 273312 57196
rect 266372 16546 266584 16574
rect 267844 16546 268424 16574
rect 269132 16546 270080 16574
rect 270512 16546 270816 16574
rect 271892 16546 272472 16574
rect 264244 3188 264296 3194
rect 264244 3130 264296 3136
rect 265348 3188 265400 3194
rect 265348 3130 265400 3136
rect 265360 480 265388 3130
rect 266556 480 266584 16546
rect 267740 3732 267792 3738
rect 267740 3674 267792 3680
rect 267752 480 267780 3674
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 16546
rect 270052 480 270080 16546
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 16546
rect 272444 480 272472 16546
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273272 354 273300 57190
rect 276020 17264 276072 17270
rect 276020 17206 276072 17212
rect 274824 5024 274876 5030
rect 274824 4966 274876 4972
rect 274836 480 274864 4966
rect 276032 480 276060 17206
rect 277412 16574 277440 84798
rect 281540 49020 281592 49026
rect 281540 48962 281592 48968
rect 280160 28280 280212 28286
rect 280160 28222 280212 28228
rect 278780 18624 278832 18630
rect 278780 18566 278832 18572
rect 278792 16574 278820 18566
rect 280172 16574 280200 28222
rect 277412 16546 278360 16574
rect 278792 16546 279096 16574
rect 280172 16546 280752 16574
rect 277124 7608 277176 7614
rect 277124 7550 277176 7556
rect 277136 480 277164 7550
rect 278332 480 278360 16546
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280724 480 280752 16546
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281552 354 281580 48962
rect 282932 16574 282960 116554
rect 289820 104168 289872 104174
rect 289820 104110 289872 104116
rect 285680 64252 285732 64258
rect 285680 64194 285732 64200
rect 284300 58676 284352 58682
rect 284300 58618 284352 58624
rect 282932 16546 283144 16574
rect 283116 480 283144 16546
rect 284312 3670 284340 58618
rect 285692 16574 285720 64194
rect 288440 62892 288492 62898
rect 288440 62834 288492 62840
rect 287060 37936 287112 37942
rect 287060 37878 287112 37884
rect 287072 16574 287100 37878
rect 288452 16574 288480 62834
rect 285692 16546 286640 16574
rect 287072 16546 287376 16574
rect 288452 16546 289032 16574
rect 284392 13116 284444 13122
rect 284392 13058 284444 13064
rect 284300 3664 284352 3670
rect 284300 3606 284352 3612
rect 284404 3482 284432 13058
rect 285036 3664 285088 3670
rect 285036 3606 285088 3612
rect 284312 3454 284432 3482
rect 284312 480 284340 3454
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285048 354 285076 3606
rect 286612 480 286640 16546
rect 285374 354 285486 480
rect 285048 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 289004 480 289032 16546
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 104110
rect 291200 60036 291252 60042
rect 291200 59978 291252 59984
rect 291212 16574 291240 59978
rect 291212 16546 291424 16574
rect 291396 480 291424 16546
rect 292592 480 292620 122266
rect 299480 120828 299532 120834
rect 299480 120770 299532 120776
rect 295340 120216 295392 120222
rect 295340 120158 295392 120164
rect 293960 68400 294012 68406
rect 293960 68342 294012 68348
rect 292672 44872 292724 44878
rect 292672 44814 292724 44820
rect 292684 16574 292712 44814
rect 293972 16574 294000 68342
rect 295352 16574 295380 120158
rect 296720 94512 296772 94518
rect 296720 94454 296772 94460
rect 296732 16574 296760 94454
rect 298100 55888 298152 55894
rect 298100 55830 298152 55836
rect 292684 16546 293264 16574
rect 293972 16546 294920 16574
rect 295352 16546 295656 16574
rect 296732 16546 297312 16574
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 294892 480 294920 16546
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 295628 354 295656 16546
rect 297284 480 297312 16546
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298112 354 298140 55830
rect 299492 3482 299520 120770
rect 305000 120760 305052 120766
rect 305000 120702 305052 120708
rect 299572 109744 299624 109750
rect 299572 109686 299624 109692
rect 299584 3670 299612 109686
rect 302240 75200 302292 75206
rect 302240 75142 302292 75148
rect 302252 16574 302280 75142
rect 303618 43480 303674 43489
rect 303618 43415 303674 43424
rect 303632 16574 303660 43415
rect 305012 16574 305040 120702
rect 302252 16546 303200 16574
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 301504 15904 301556 15910
rect 301504 15846 301556 15852
rect 299572 3664 299624 3670
rect 299572 3606 299624 3612
rect 300768 3664 300820 3670
rect 300768 3606 300820 3612
rect 299492 3454 299704 3482
rect 299676 480 299704 3454
rect 300780 480 300808 3606
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 15846
rect 303172 480 303200 16546
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306392 354 306420 124170
rect 325700 122256 325752 122262
rect 325700 122198 325752 122204
rect 313280 121644 313332 121650
rect 313280 121586 313332 121592
rect 307852 100020 307904 100026
rect 307852 99962 307904 99968
rect 307024 61396 307076 61402
rect 307024 61338 307076 61344
rect 307036 3398 307064 61338
rect 307864 16574 307892 99962
rect 309138 57216 309194 57225
rect 309138 57151 309194 57160
rect 309152 16574 309180 57151
rect 310520 42084 310572 42090
rect 310520 42026 310572 42032
rect 310532 16574 310560 42026
rect 311164 33788 311216 33794
rect 311164 33730 311216 33736
rect 307864 16546 307984 16574
rect 309152 16546 309824 16574
rect 310532 16546 311112 16574
rect 307024 3392 307076 3398
rect 307024 3334 307076 3340
rect 307956 480 307984 16546
rect 309048 3392 309100 3398
rect 309048 3334 309100 3340
rect 309060 480 309088 3334
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 16546
rect 311084 3482 311112 16546
rect 311176 3670 311204 33730
rect 313292 16574 313320 121586
rect 314660 115252 314712 115258
rect 314660 115194 314712 115200
rect 313292 16546 313872 16574
rect 311164 3664 311216 3670
rect 311164 3606 311216 3612
rect 312636 3664 312688 3670
rect 312636 3606 312688 3612
rect 311084 3454 311480 3482
rect 311452 480 311480 3454
rect 312648 480 312676 3606
rect 313844 480 313872 16546
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314672 354 314700 115194
rect 317420 113824 317472 113830
rect 317420 113766 317472 113772
rect 316040 87644 316092 87650
rect 316040 87586 316092 87592
rect 316052 3398 316080 87586
rect 316132 22772 316184 22778
rect 316132 22714 316184 22720
rect 316144 16574 316172 22714
rect 317432 16574 317460 113766
rect 324320 95260 324372 95266
rect 324320 95202 324372 95208
rect 320180 64184 320232 64190
rect 320180 64126 320232 64132
rect 320192 16574 320220 64126
rect 322940 31068 322992 31074
rect 322940 31010 322992 31016
rect 316144 16546 316264 16574
rect 317432 16546 318104 16574
rect 320192 16546 320496 16574
rect 316040 3392 316092 3398
rect 316040 3334 316092 3340
rect 316236 480 316264 16546
rect 317328 3392 317380 3398
rect 317328 3334 317380 3340
rect 317340 480 317368 3334
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319720 3596 319772 3602
rect 319720 3538 319772 3544
rect 319732 480 319760 3538
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322112 4956 322164 4962
rect 322112 4898 322164 4904
rect 322124 480 322152 4898
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 31010
rect 324332 3602 324360 95202
rect 325712 16574 325740 122198
rect 580356 120148 580408 120154
rect 580356 120090 580408 120096
rect 349160 118720 349212 118726
rect 349160 118662 349212 118668
rect 336740 108316 336792 108322
rect 336740 108258 336792 108264
rect 329840 89004 329892 89010
rect 329840 88946 329892 88952
rect 327080 62824 327132 62830
rect 327080 62766 327132 62772
rect 327092 16574 327120 62766
rect 328458 58576 328514 58585
rect 328458 58511 328514 58520
rect 328472 16574 328500 58511
rect 329852 16574 329880 88946
rect 332600 84244 332652 84250
rect 332600 84186 332652 84192
rect 331220 83496 331272 83502
rect 331220 83438 331272 83444
rect 325712 16546 326384 16574
rect 327092 16546 328040 16574
rect 328472 16546 328776 16574
rect 329852 16546 330432 16574
rect 324412 4888 324464 4894
rect 324412 4830 324464 4836
rect 324320 3596 324372 3602
rect 324320 3538 324372 3544
rect 324424 480 324452 4830
rect 325608 3596 325660 3602
rect 325608 3538 325660 3544
rect 325620 480 325648 3538
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 16546
rect 328012 480 328040 16546
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 328748 354 328776 16546
rect 330404 480 330432 16546
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 83438
rect 332612 3482 332640 84186
rect 333980 51740 334032 51746
rect 333980 51682 334032 51688
rect 332690 19952 332746 19961
rect 332690 19887 332746 19896
rect 332704 3602 332732 19887
rect 333992 16574 334020 51682
rect 335358 40624 335414 40633
rect 335358 40559 335414 40568
rect 335372 16574 335400 40559
rect 336752 16574 336780 108258
rect 347780 106956 347832 106962
rect 347780 106898 347832 106904
rect 346400 90364 346452 90370
rect 346400 90306 346452 90312
rect 339500 74588 339552 74594
rect 339500 74530 339552 74536
rect 338118 54496 338174 54505
rect 338118 54431 338174 54440
rect 338132 16574 338160 54431
rect 333992 16546 334664 16574
rect 335372 16546 336320 16574
rect 336752 16546 337056 16574
rect 338132 16546 338712 16574
rect 332692 3596 332744 3602
rect 332692 3538 332744 3544
rect 333888 3596 333940 3602
rect 333888 3538 333940 3544
rect 332612 3454 332732 3482
rect 332704 480 332732 3454
rect 333900 480 333928 3538
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 336292 480 336320 16546
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338684 480 338712 16546
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 74530
rect 340970 53136 341026 53145
rect 340970 53071 341026 53080
rect 340984 3534 341012 53071
rect 345020 47592 345072 47598
rect 345020 47534 345072 47540
rect 345032 16574 345060 47534
rect 346412 16574 346440 90306
rect 347792 16574 347820 106898
rect 345032 16546 345336 16574
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 343364 4820 343416 4826
rect 343364 4762 343416 4768
rect 340972 3528 341024 3534
rect 340972 3470 341024 3476
rect 342168 3528 342220 3534
rect 342168 3470 342220 3476
rect 340972 3392 341024 3398
rect 340972 3334 341024 3340
rect 340984 480 341012 3334
rect 342180 480 342208 3470
rect 343376 480 343404 4762
rect 344560 3596 344612 3602
rect 344560 3538 344612 3544
rect 344572 480 344600 3538
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 346964 480 346992 16546
rect 348068 480 348096 16546
rect 349172 3534 349200 118662
rect 580264 117972 580316 117978
rect 580264 117914 580316 117920
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580184 99414 580212 99447
rect 580172 99408 580224 99414
rect 580172 99350 580224 99356
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580184 85610 580212 86119
rect 580172 85604 580224 85610
rect 580172 85546 580224 85552
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580184 71806 580212 72927
rect 580172 71800 580224 71806
rect 580172 71742 580224 71748
rect 350540 68332 350592 68338
rect 350540 68274 350592 68280
rect 349252 66904 349304 66910
rect 349252 66846 349304 66852
rect 349160 3528 349212 3534
rect 349160 3470 349212 3476
rect 349264 480 349292 66846
rect 350552 16574 350580 68274
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 580276 19825 580304 117914
rect 580368 112849 580396 120090
rect 580354 112840 580410 112849
rect 580354 112775 580410 112784
rect 580262 19816 580318 19825
rect 580262 19751 580318 19760
rect 350552 16546 351224 16574
rect 350448 3528 350500 3534
rect 350448 3470 350500 3476
rect 350460 480 350488 3470
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3054 501744 3110 501800
rect 2778 475632 2834 475688
rect 3238 462576 3294 462632
rect 3146 449520 3202 449576
rect 3422 423544 3478 423600
rect 3422 410488 3478 410544
rect 3330 345344 3386 345400
rect 3330 319232 3386 319288
rect 3330 293120 3386 293176
rect 3514 397468 3516 397488
rect 3516 397468 3568 397488
rect 3568 397468 3570 397488
rect 3514 397432 3570 397468
rect 3606 371320 3662 371376
rect 3514 358400 3570 358456
rect 3422 267144 3478 267200
rect 3146 254088 3202 254144
rect 3054 241032 3110 241088
rect 3330 214920 3386 214976
rect 3698 306176 3754 306232
rect 3514 206216 3570 206272
rect 3422 201864 3478 201920
rect 54482 198600 54538 198656
rect 3422 188808 3478 188864
rect 3422 162832 3478 162888
rect 2962 149776 3018 149832
rect 3514 136720 3570 136776
rect 3422 110608 3478 110664
rect 3422 84632 3478 84688
rect 2870 71576 2926 71632
rect 2778 45500 2780 45520
rect 2780 45500 2832 45520
rect 2832 45500 2834 45520
rect 2778 45464 2834 45500
rect 2870 32408 2926 32464
rect 3606 97552 3662 97608
rect 3514 58520 3570 58576
rect 64694 251368 64750 251424
rect 65338 210160 65394 210216
rect 65430 200232 65486 200288
rect 65982 251504 66038 251560
rect 66074 112104 66130 112160
rect 66902 223760 66958 223816
rect 66902 197920 66958 197976
rect 67638 247716 67694 247752
rect 67638 247696 67640 247716
rect 67640 247696 67692 247716
rect 67692 247696 67694 247716
rect 67546 245520 67602 245576
rect 67454 241576 67510 241632
rect 67638 244316 67694 244352
rect 67638 244296 67640 244316
rect 67640 244296 67692 244316
rect 67692 244296 67694 244316
rect 68282 245520 68338 245576
rect 68374 240932 68376 240952
rect 68376 240932 68428 240952
rect 68428 240932 68430 240952
rect 68374 240896 68430 240932
rect 66994 104080 67050 104136
rect 66810 83544 66866 83600
rect 67638 230560 67694 230616
rect 67730 229336 67786 229392
rect 68374 236816 68430 236872
rect 68558 247696 68614 247752
rect 68374 232056 68430 232112
rect 68466 227976 68522 228032
rect 67822 225800 67878 225856
rect 68190 225800 68246 225856
rect 68006 221040 68062 221096
rect 67270 101360 67326 101416
rect 68190 219000 68246 219056
rect 68466 218320 68522 218376
rect 68374 216960 68430 217016
rect 67638 216280 67694 216336
rect 68374 214920 68430 214976
rect 67638 214376 67694 214432
rect 68190 214376 68246 214432
rect 67914 213560 67970 213616
rect 67730 206216 67786 206272
rect 67638 202680 67694 202736
rect 67822 205572 67824 205592
rect 67824 205572 67876 205592
rect 67876 205572 67878 205592
rect 67822 205536 67878 205572
rect 68098 204720 68154 204776
rect 68374 201184 68430 201240
rect 68742 249736 68798 249792
rect 68650 243616 68706 243672
rect 68834 248240 68890 248296
rect 68834 237496 68890 237552
rect 68742 232620 68798 232656
rect 68742 232600 68744 232620
rect 68744 232600 68796 232620
rect 68796 232600 68798 232620
rect 68650 230016 68706 230072
rect 69110 246200 69166 246256
rect 69018 234096 69074 234152
rect 68926 227296 68982 227352
rect 68742 225292 68744 225312
rect 68744 225292 68796 225312
rect 68796 225292 68798 225312
rect 68742 225256 68798 225292
rect 69018 225256 69074 225312
rect 68650 223080 68706 223136
rect 68926 220360 68982 220416
rect 68650 201320 68706 201376
rect 68190 186632 68246 186688
rect 67730 180920 67786 180976
rect 67546 105440 67602 105496
rect 67638 104796 67640 104816
rect 67640 104796 67692 104816
rect 67692 104796 67694 104816
rect 67638 104760 67694 104796
rect 67638 102720 67694 102776
rect 67638 100700 67694 100736
rect 67638 100680 67640 100700
rect 67640 100680 67692 100700
rect 67692 100680 67694 100700
rect 67638 98640 67694 98696
rect 67638 97824 67694 97880
rect 67638 95920 67694 95976
rect 67638 93200 67694 93256
rect 67638 91160 67694 91216
rect 67638 84360 67694 84416
rect 67638 78784 67694 78840
rect 67638 78240 67694 78296
rect 67638 77596 67640 77616
rect 67640 77596 67692 77616
rect 67692 77596 67694 77616
rect 67638 77560 67694 77596
rect 67914 87760 67970 87816
rect 67914 85720 67970 85776
rect 67822 80824 67878 80880
rect 67730 75792 67786 75848
rect 68098 91840 68154 91896
rect 68098 86980 68100 87000
rect 68100 86980 68152 87000
rect 68152 86980 68154 87000
rect 68098 86944 68154 86980
rect 68834 208120 68890 208176
rect 68926 204856 68982 204912
rect 68926 177284 68928 177304
rect 68928 177284 68980 177304
rect 68980 177284 68982 177304
rect 68926 177248 68982 177284
rect 68558 106800 68614 106856
rect 68282 100000 68338 100056
rect 68558 88984 68614 89040
rect 68466 88476 68468 88496
rect 68468 88476 68520 88496
rect 68520 88476 68522 88496
rect 68466 88440 68522 88476
rect 68190 80824 68246 80880
rect 68006 78784 68062 78840
rect 68282 71984 68338 72040
rect 68466 81504 68522 81560
rect 68834 117272 68890 117328
rect 68834 116048 68890 116104
rect 68834 107480 68890 107536
rect 68926 94560 68982 94616
rect 71962 251776 72018 251832
rect 73066 251776 73122 251832
rect 78402 249872 78458 249928
rect 84198 251504 84254 251560
rect 82266 250008 82322 250064
rect 84842 251368 84898 251424
rect 88706 250144 88762 250200
rect 94686 251640 94742 251696
rect 95146 250416 95202 250472
rect 103426 251096 103482 251152
rect 106094 251912 106150 251968
rect 112166 249736 112222 249792
rect 119158 252864 119214 252920
rect 116398 251232 116454 251288
rect 118698 251368 118754 251424
rect 119250 251640 119306 251696
rect 119342 249872 119398 249928
rect 69478 243500 69534 243536
rect 69478 243480 69480 243500
rect 69480 243480 69532 243500
rect 69532 243480 69534 243500
rect 69386 236136 69442 236192
rect 69294 234776 69350 234832
rect 119894 251776 119950 251832
rect 119342 230968 119398 231024
rect 69478 221720 69534 221776
rect 69386 211520 69442 211576
rect 69294 200640 69350 200696
rect 69662 211928 69718 211984
rect 119342 219544 119398 219600
rect 119526 218476 119582 218512
rect 119526 218456 119528 218476
rect 119528 218456 119580 218476
rect 119580 218456 119582 218476
rect 70674 200232 70730 200288
rect 69386 175924 69388 175944
rect 69388 175924 69440 175944
rect 69440 175924 69442 175944
rect 69386 175888 69442 175924
rect 69110 105984 69166 106040
rect 69018 88984 69074 89040
rect 68834 86264 68890 86320
rect 68926 75792 68982 75848
rect 68926 74840 68982 74896
rect 68650 71304 68706 71360
rect 68466 67224 68522 67280
rect 68282 65728 68338 65784
rect 68834 74024 68890 74080
rect 3514 19352 3570 19408
rect 3422 6432 3478 6488
rect 69202 95240 69258 95296
rect 69570 99320 69626 99376
rect 69846 111560 69902 111616
rect 70306 109928 70362 109984
rect 70214 108568 70270 108624
rect 69662 97280 69718 97336
rect 69478 93880 69534 93936
rect 69386 90480 69442 90536
rect 69294 86944 69350 87000
rect 69294 82184 69350 82240
rect 69202 69672 69258 69728
rect 69754 80144 69810 80200
rect 69386 79464 69442 79520
rect 69478 76744 69534 76800
rect 69570 73208 69626 73264
rect 69570 72664 69626 72720
rect 69662 70624 69718 70680
rect 69570 64776 69626 64832
rect 69846 71304 69902 71360
rect 70490 199824 70546 199880
rect 72606 198736 72662 198792
rect 82082 199300 82138 199336
rect 82082 199280 82084 199300
rect 82084 199280 82136 199300
rect 82136 199280 82138 199300
rect 84934 199316 84936 199336
rect 84936 199316 84988 199336
rect 84988 199316 84990 199336
rect 84934 199280 84990 199316
rect 74538 168952 74594 169008
rect 93858 198056 93914 198112
rect 103426 198464 103482 198520
rect 76470 117952 76526 118008
rect 73250 116184 73306 116240
rect 74998 112104 75054 112160
rect 74998 111832 75054 111888
rect 76470 116456 76526 116512
rect 106186 77152 106242 77208
rect 106186 76472 106242 76528
rect 106186 74976 106242 75032
rect 70306 69944 70362 70000
rect 70398 67904 70454 67960
rect 74538 68176 74594 68232
rect 77758 68720 77814 68776
rect 78402 65864 78458 65920
rect 79690 68312 79746 68368
rect 84198 68448 84254 68504
rect 89350 68856 89406 68912
rect 88062 67088 88118 67144
rect 95146 68584 95202 68640
rect 100942 67360 100998 67416
rect 106186 70352 106242 70408
rect 107474 198600 107530 198656
rect 106370 108432 106426 108488
rect 103518 66136 103574 66192
rect 106278 66000 106334 66056
rect 106462 104760 106518 104816
rect 106462 102312 106518 102368
rect 106554 97824 106610 97880
rect 107014 168952 107070 169008
rect 107658 108996 107714 109032
rect 107658 108976 107660 108996
rect 107660 108976 107712 108996
rect 107712 108976 107714 108996
rect 108026 108432 108082 108488
rect 108026 104796 108028 104816
rect 108028 104796 108080 104816
rect 108080 104796 108082 104816
rect 108026 104760 108082 104796
rect 107658 98912 107714 98968
rect 107750 97824 107806 97880
rect 107658 97552 107714 97608
rect 107750 96464 107806 96520
rect 107658 96192 107714 96248
rect 107842 95512 107898 95568
rect 107658 94832 107714 94888
rect 107658 94152 107714 94208
rect 107658 93472 107714 93528
rect 107750 92792 107806 92848
rect 107750 91432 107806 91488
rect 107658 90072 107714 90128
rect 108026 90752 108082 90808
rect 107014 66000 107070 66056
rect 107566 65728 107622 65784
rect 107750 79872 107806 79928
rect 107750 77832 107806 77888
rect 107750 77188 107752 77208
rect 107752 77188 107804 77208
rect 107804 77188 107806 77208
rect 107750 77152 107806 77188
rect 107750 75948 107806 75984
rect 107750 75928 107752 75948
rect 107752 75928 107804 75948
rect 107804 75928 107806 75948
rect 107842 75792 107898 75848
rect 107750 75148 107752 75168
rect 107752 75148 107804 75168
rect 107804 75148 107806 75168
rect 107750 75112 107806 75148
rect 107750 74468 107752 74488
rect 107752 74468 107804 74488
rect 107804 74468 107806 74488
rect 107750 74432 107806 74468
rect 107842 73072 107898 73128
rect 107750 72392 107806 72448
rect 108210 104352 108266 104408
rect 108210 102312 108266 102368
rect 108210 84632 108266 84688
rect 108578 196560 108634 196616
rect 108854 196696 108910 196752
rect 108578 109792 108634 109848
rect 108762 100952 108818 101008
rect 108762 99592 108818 99648
rect 108670 89392 108726 89448
rect 108578 88712 108634 88768
rect 108486 87352 108542 87408
rect 108578 85992 108634 86048
rect 108946 111152 109002 111208
rect 108946 110372 108948 110392
rect 108948 110372 109000 110392
rect 109000 110372 109002 110392
rect 108946 110336 109002 110372
rect 108946 107072 109002 107128
rect 108946 106392 109002 106448
rect 108946 105712 109002 105768
rect 108946 102992 109002 103048
rect 108946 101632 109002 101688
rect 108946 100272 109002 100328
rect 108946 88032 109002 88088
rect 108946 86672 109002 86728
rect 108946 83952 109002 84008
rect 108946 82592 109002 82648
rect 108854 81912 108910 81968
rect 108854 81268 108856 81288
rect 108856 81268 108908 81288
rect 108908 81268 108910 81288
rect 108854 81232 108910 81268
rect 108946 80552 109002 80608
rect 108670 79228 108672 79248
rect 108672 79228 108724 79248
rect 108724 79228 108726 79248
rect 108670 79192 108726 79228
rect 109222 83272 109278 83328
rect 109774 87488 109830 87544
rect 111522 123392 111578 123448
rect 112994 192480 113050 192536
rect 112902 175888 112958 175944
rect 113086 73752 113142 73808
rect 113086 71032 113142 71088
rect 111246 68176 111302 68232
rect 113546 69400 113602 69456
rect 113822 69264 113878 69320
rect 113362 68584 113418 68640
rect 114650 68448 114706 68504
rect 116582 71032 116638 71088
rect 115938 68856 115994 68912
rect 115846 68448 115902 68504
rect 117042 124480 117098 124536
rect 119710 199416 119766 199472
rect 119342 165552 119398 165608
rect 119250 125432 119306 125488
rect 119710 125296 119766 125352
rect 120170 219816 120226 219872
rect 120170 217640 120226 217696
rect 120078 203360 120134 203416
rect 120446 220360 120502 220416
rect 120354 201320 120410 201376
rect 121458 248240 121514 248296
rect 121458 246880 121514 246936
rect 121458 244296 121514 244352
rect 121642 244840 121698 244896
rect 121458 242120 121514 242176
rect 121550 241596 121606 241632
rect 121550 241576 121552 241596
rect 121552 241576 121604 241596
rect 121604 241576 121606 241596
rect 121458 238040 121514 238096
rect 120722 208120 120778 208176
rect 120630 166912 120686 166968
rect 119986 95240 120042 95296
rect 121458 230696 121514 230752
rect 121458 229200 121514 229256
rect 121458 224576 121514 224632
rect 121550 222536 121606 222592
rect 121458 221856 121514 221912
rect 121458 215736 121514 215792
rect 121458 214920 121514 214976
rect 121458 212200 121514 212256
rect 121550 210976 121606 211032
rect 121550 206760 121606 206816
rect 121550 206080 121606 206136
rect 121826 239536 121882 239592
rect 121826 237360 121882 237416
rect 121734 232736 121790 232792
rect 121734 213016 121790 213072
rect 122010 246200 122066 246256
rect 122378 248920 122434 248976
rect 122654 245792 122710 245848
rect 122286 242972 122288 242992
rect 122288 242972 122340 242992
rect 122340 242972 122342 242992
rect 122286 242936 122342 242972
rect 121918 222536 121974 222592
rect 122010 216960 122066 217016
rect 121918 213560 121974 213616
rect 122286 235320 122342 235376
rect 122470 234660 122526 234696
rect 122470 234640 122472 234660
rect 122472 234640 122524 234660
rect 122524 234640 122526 234660
rect 122470 233300 122526 233336
rect 122470 233280 122472 233300
rect 122472 233280 122524 233300
rect 122524 233280 122526 233300
rect 122194 223760 122250 223816
rect 121734 205400 121790 205456
rect 121826 202000 121882 202056
rect 117226 68856 117282 68912
rect 117226 68448 117282 68504
rect 116674 68312 116730 68368
rect 115846 68040 115902 68096
rect 113914 65864 113970 65920
rect 122470 225800 122526 225856
rect 122378 208800 122434 208856
rect 122562 205400 122618 205456
rect 122562 204040 122618 204096
rect 122562 201320 122618 201376
rect 122746 236020 122802 236056
rect 122746 236000 122748 236020
rect 122748 236000 122800 236020
rect 122800 236000 122802 236020
rect 123574 252728 123630 252784
rect 123758 252592 123814 252648
rect 122838 198464 122894 198520
rect 122194 122848 122250 122904
rect 131118 251252 131174 251288
rect 131118 251232 131120 251252
rect 131120 251232 131172 251252
rect 131172 251232 131174 251252
rect 131118 121388 131120 121408
rect 131120 121388 131172 121408
rect 131172 121388 131174 121408
rect 131118 121352 131174 121388
rect 133142 247560 133198 247616
rect 131854 121352 131910 121408
rect 133786 247560 133842 247616
rect 140778 232464 140834 232520
rect 140778 113736 140834 113792
rect 141422 113736 141478 113792
rect 141514 67360 141570 67416
rect 143446 114028 143502 114064
rect 143446 114008 143448 114028
rect 143448 114008 143500 114028
rect 143500 114008 143502 114028
rect 145562 97960 145618 98016
rect 152462 250552 152518 250608
rect 150438 112240 150494 112296
rect 153014 113892 153070 113928
rect 153014 113872 153016 113892
rect 153016 113872 153068 113892
rect 153068 113872 153070 113892
rect 153106 73888 153162 73944
rect 156786 165552 156842 165608
rect 162030 112104 162086 112160
rect 162674 96464 162730 96520
rect 163410 68856 163466 68912
rect 164882 168000 164938 168056
rect 164146 122032 164202 122088
rect 164698 112240 164754 112296
rect 164698 111832 164754 111888
rect 165434 169496 165490 169552
rect 164054 68856 164110 68912
rect 163870 68720 163926 68776
rect 163410 67904 163466 67960
rect 166538 167728 166594 167784
rect 165986 122168 166042 122224
rect 165342 67496 165398 67552
rect 165526 67496 165582 67552
rect 165526 67088 165582 67144
rect 166538 121896 166594 121952
rect 166262 68040 166318 68096
rect 166998 229200 167054 229256
rect 166906 119584 166962 119640
rect 167090 227840 167146 227896
rect 167090 225800 167146 225856
rect 167090 224440 167146 224496
rect 167090 223080 167146 223136
rect 167090 219000 167146 219056
rect 167090 217640 167146 217696
rect 167090 216280 167146 216336
rect 167182 214920 167238 214976
rect 167090 214240 167146 214296
rect 167090 211540 167146 211576
rect 167090 211520 167092 211540
rect 167092 211520 167144 211540
rect 167144 211520 167146 211540
rect 167550 227160 167606 227216
rect 167458 221040 167514 221096
rect 167366 211520 167422 211576
rect 167090 210860 167146 210896
rect 167090 210840 167092 210860
rect 167092 210840 167144 210860
rect 167144 210840 167146 210860
rect 167274 210840 167330 210896
rect 167826 222400 167882 222456
rect 167734 219680 167790 219736
rect 167642 212880 167698 212936
rect 167090 208120 167146 208176
rect 167090 206760 167146 206816
rect 167090 206080 167146 206136
rect 167090 201320 167146 201376
rect 167366 206080 167422 206136
rect 167274 203360 167330 203416
rect 167458 202680 167514 202736
rect 167366 199960 167422 200016
rect 167366 197920 167422 197976
rect 167366 196596 167368 196616
rect 167368 196596 167420 196616
rect 167420 196596 167422 196616
rect 167366 196560 167422 196596
rect 167366 191800 167422 191856
rect 167366 189760 167422 189816
rect 167366 186380 167422 186416
rect 167366 186360 167368 186380
rect 167368 186360 167420 186380
rect 167420 186360 167422 186380
rect 167366 185000 167422 185056
rect 167366 183640 167422 183696
rect 167366 182280 167422 182336
rect 167458 180240 167514 180296
rect 167458 176840 167514 176896
rect 168194 209480 168250 209536
rect 168286 206760 168342 206816
rect 168930 198192 168986 198248
rect 168194 195200 168250 195256
rect 168286 193160 168342 193216
rect 168102 190440 168158 190496
rect 168286 185000 168342 185056
rect 168194 180240 168250 180296
rect 168102 175480 168158 175536
rect 168102 172080 168158 172136
rect 168102 170720 168158 170776
rect 167274 118768 167330 118824
rect 167090 118224 167146 118280
rect 166998 117544 167054 117600
rect 166998 115504 167054 115560
rect 167182 114860 167184 114880
rect 167184 114860 167236 114880
rect 167236 114860 167238 114880
rect 167182 114824 167238 114860
rect 166998 112104 167054 112160
rect 166906 111832 166962 111888
rect 166998 110200 167054 110256
rect 167090 109520 167146 109576
rect 166998 107480 167054 107536
rect 166998 106664 167054 106720
rect 166998 103436 167000 103456
rect 167000 103436 167052 103456
rect 167052 103436 167054 103456
rect 166998 103400 167054 103436
rect 166998 102076 167000 102096
rect 167000 102076 167052 102096
rect 167052 102076 167054 102096
rect 166998 102040 167054 102076
rect 167458 100700 167514 100736
rect 167458 100680 167460 100700
rect 167460 100680 167512 100700
rect 167512 100680 167514 100700
rect 167090 100000 167146 100056
rect 167550 98640 167606 98696
rect 167182 97860 167184 97880
rect 167184 97860 167236 97880
rect 167236 97860 167238 97880
rect 167182 97824 167238 97860
rect 166998 94560 167054 94616
rect 166906 93200 166962 93256
rect 167274 92520 167330 92576
rect 166998 89800 167054 89856
rect 166998 88984 167054 89040
rect 167182 88440 167238 88496
rect 167090 87760 167146 87816
rect 166998 85604 167054 85640
rect 166998 85584 167000 85604
rect 167000 85584 167052 85604
rect 167052 85584 167054 85604
rect 167090 84360 167146 84416
rect 166998 83000 167054 83056
rect 166998 81504 167054 81560
rect 166998 80280 167054 80336
rect 166998 78804 167054 78840
rect 166998 78784 167000 78804
rect 167000 78784 167052 78804
rect 167052 78784 167054 78804
rect 166814 69536 166870 69592
rect 166354 67224 166410 67280
rect 167090 74704 167146 74760
rect 167090 74024 167146 74080
rect 167182 73344 167238 73400
rect 167090 71984 167146 72040
rect 167918 105440 167974 105496
rect 167734 93880 167790 93936
rect 167734 91160 167790 91216
rect 167642 90480 167698 90536
rect 167918 92520 167974 92576
rect 167642 79464 167698 79520
rect 167458 70352 167514 70408
rect 167734 78104 167790 78160
rect 168010 71304 168066 71360
rect 168746 173440 168802 173496
rect 169114 173440 169170 173496
rect 168930 168136 168986 168192
rect 168746 167864 168802 167920
rect 168654 121760 168710 121816
rect 168470 120536 168526 120592
rect 168378 120264 168434 120320
rect 168930 116048 168986 116104
rect 168930 108840 168986 108896
rect 169206 118224 169262 118280
rect 169114 116084 169116 116104
rect 169116 116084 169168 116104
rect 169168 116084 169170 116104
rect 169114 116048 169170 116084
rect 169298 114144 169354 114200
rect 169114 106120 169170 106176
rect 169022 104760 169078 104816
rect 169206 104080 169262 104136
rect 169022 100680 169078 100736
rect 168930 97824 168986 97880
rect 168838 95240 168894 95296
rect 168286 79464 168342 79520
rect 168286 77424 168342 77480
rect 168194 76880 168250 76936
rect 168102 70624 168158 70680
rect 169114 98640 169170 98696
rect 169390 112784 169446 112840
rect 169574 190440 169630 190496
rect 169942 194520 169998 194576
rect 171230 230560 171286 230616
rect 178038 250416 178094 250472
rect 182178 249736 182234 249792
rect 182822 249736 182878 249792
rect 183558 233144 183614 233200
rect 187054 247968 187110 248024
rect 184202 233144 184258 233200
rect 229282 228792 229338 228848
rect 229282 227704 229338 227760
rect 229282 209208 229338 209264
rect 170126 204992 170182 205048
rect 229466 228792 229522 228848
rect 229834 228928 229890 228984
rect 229650 226616 229706 226672
rect 229558 212472 229614 212528
rect 229374 202952 229430 203008
rect 169850 188944 169906 189000
rect 169666 179288 169722 179344
rect 229374 196152 229430 196208
rect 170310 169632 170366 169688
rect 175186 168952 175242 169008
rect 170954 168272 171010 168328
rect 182914 167864 182970 167920
rect 184938 168272 184994 168328
rect 193218 168000 193274 168056
rect 198370 169496 198426 169552
rect 199658 168272 199714 168328
rect 169942 121624 169998 121680
rect 175186 120128 175242 120184
rect 178406 121896 178462 121952
rect 180982 121624 181038 121680
rect 180338 120536 180394 120592
rect 182270 120400 182326 120456
rect 186778 122032 186834 122088
rect 191286 122168 191342 122224
rect 188710 120264 188766 120320
rect 192574 121760 192630 121816
rect 193126 121352 193182 121408
rect 193218 120672 193274 120728
rect 170678 119312 170734 119368
rect 169574 116048 169630 116104
rect 169482 110744 169538 110800
rect 169390 109520 169446 109576
rect 169482 100000 169538 100056
rect 200118 119312 200174 119368
rect 200118 113056 200174 113112
rect 200302 113056 200358 113112
rect 169850 106120 169906 106176
rect 169758 88440 169814 88496
rect 200118 104352 200174 104408
rect 200118 98232 200174 98288
rect 200394 110472 200450 110528
rect 200302 108432 200358 108488
rect 200210 95512 200266 95568
rect 201406 95512 201462 95568
rect 200210 94832 200266 94888
rect 200302 92792 200358 92848
rect 200118 85992 200174 86048
rect 198738 70624 198794 70680
rect 170034 70352 170090 70408
rect 171322 68856 171378 68912
rect 171874 68856 171930 68912
rect 174542 68176 174598 68232
rect 173254 66000 173310 66056
rect 177302 68720 177358 68776
rect 177762 68720 177818 68776
rect 179694 68312 179750 68368
rect 180062 68312 180118 68368
rect 178406 65864 178462 65920
rect 189078 68856 189134 68912
rect 189078 68448 189134 68504
rect 188710 67496 188766 67552
rect 190366 68856 190422 68912
rect 192574 68584 192630 68640
rect 199382 69808 199438 69864
rect 200118 85584 200174 85640
rect 200210 71848 200266 71904
rect 201590 105712 201646 105768
rect 201958 118632 202014 118688
rect 201958 117972 202014 118008
rect 201958 117952 201960 117972
rect 201960 117952 202012 117972
rect 202012 117952 202014 117972
rect 201958 115252 202014 115288
rect 201958 115232 201960 115252
rect 201960 115232 202012 115252
rect 202012 115232 202014 115252
rect 201866 111832 201922 111888
rect 202142 117272 202198 117328
rect 202418 115776 202474 115832
rect 202326 114416 202382 114472
rect 202050 111152 202106 111208
rect 201866 109812 201922 109848
rect 201866 109792 201868 109812
rect 201868 109792 201920 109812
rect 201920 109792 201922 109812
rect 202786 109112 202842 109168
rect 202786 107072 202842 107128
rect 202234 106392 202290 106448
rect 201774 105032 201830 105088
rect 201866 103672 201922 103728
rect 201682 102992 201738 103048
rect 201590 100272 201646 100328
rect 201590 98912 201646 98968
rect 201866 101632 201922 101688
rect 201498 82864 201554 82920
rect 200670 77288 200726 77344
rect 200486 75112 200542 75168
rect 200578 73208 200634 73264
rect 200210 67360 200266 67416
rect 201314 76472 201370 76528
rect 200946 74704 201002 74760
rect 200854 73752 200910 73808
rect 200762 72392 200818 72448
rect 202786 99592 202842 99648
rect 201958 97552 202014 97608
rect 201774 90788 201776 90808
rect 201776 90788 201828 90808
rect 201828 90788 201830 90808
rect 201774 90752 201830 90788
rect 201774 90092 201830 90128
rect 201774 90072 201776 90092
rect 201776 90072 201828 90092
rect 201828 90072 201830 90092
rect 202142 96464 202198 96520
rect 202418 96192 202474 96248
rect 202050 92112 202106 92168
rect 202142 89392 202198 89448
rect 202050 80552 202106 80608
rect 201958 73752 202014 73808
rect 201958 71168 202014 71224
rect 202050 70488 202106 70544
rect 202234 81912 202290 81968
rect 202786 94152 202842 94208
rect 202510 88712 202566 88768
rect 202510 88032 202566 88088
rect 202510 86672 202566 86728
rect 202694 84804 202696 84824
rect 202696 84804 202748 84824
rect 202748 84804 202750 84824
rect 202694 84768 202750 84804
rect 202694 84244 202750 84280
rect 202694 84224 202696 84244
rect 202696 84224 202748 84244
rect 202748 84224 202750 84244
rect 202510 80144 202566 80200
rect 202786 79192 202842 79248
rect 202786 78684 202788 78704
rect 202788 78684 202840 78704
rect 202840 78684 202842 78704
rect 202786 78648 202842 78684
rect 202510 69672 202566 69728
rect 200854 66136 200910 66192
rect 203154 83272 203210 83328
rect 204442 122848 204498 122904
rect 218334 168156 218390 168192
rect 218334 168136 218336 168156
rect 218336 168136 218388 168156
rect 218388 168136 218390 168156
rect 221554 169632 221610 169688
rect 226062 167728 226118 167784
rect 229282 169496 229338 169552
rect 229466 195336 229522 195392
rect 229558 192752 229614 192808
rect 230294 227160 230350 227216
rect 230202 225800 230258 225856
rect 230110 221040 230166 221096
rect 230018 219000 230074 219056
rect 230570 212880 230626 212936
rect 230570 212200 230626 212256
rect 230478 210840 230534 210896
rect 230386 209480 230442 209536
rect 230018 207440 230074 207496
rect 229926 204040 229982 204096
rect 229742 181056 229798 181112
rect 230754 214240 230810 214296
rect 230662 206080 230718 206136
rect 230938 222400 230994 222456
rect 231306 223760 231362 223816
rect 231398 220360 231454 220416
rect 231214 216960 231270 217016
rect 231122 215600 231178 215656
rect 231030 174800 231086 174856
rect 231858 185000 231914 185056
rect 231858 179560 231914 179616
rect 231766 171828 231822 171864
rect 231766 171808 231768 171828
rect 231768 171808 231820 171828
rect 231820 171808 231822 171828
rect 231674 171128 231730 171184
rect 232686 225120 232742 225176
rect 232686 217948 232688 217968
rect 232688 217948 232740 217968
rect 232740 217948 232742 217968
rect 232686 217912 232742 217948
rect 232686 206080 232742 206136
rect 233146 204720 233202 204776
rect 232686 204040 232742 204096
rect 232686 202680 232742 202736
rect 232594 200640 232650 200696
rect 232686 199280 232742 199336
rect 232594 197920 232650 197976
rect 232410 194520 232466 194576
rect 232318 192480 232374 192536
rect 232226 189760 232282 189816
rect 232134 184320 232190 184376
rect 232410 182960 232466 183016
rect 232226 180240 232282 180296
rect 232042 178200 232098 178256
rect 231950 176160 232006 176216
rect 232042 173440 232098 173496
rect 232502 176840 232558 176896
rect 233146 191140 233202 191176
rect 233146 191120 233148 191140
rect 233148 191120 233200 191140
rect 233200 191120 233202 191140
rect 232778 188400 232834 188456
rect 233146 187720 233202 187776
rect 233146 186360 233202 186416
rect 233054 174800 233110 174856
rect 233330 201320 233386 201376
rect 233330 166912 233386 166968
rect 233882 170040 233938 170096
rect 233606 165552 233662 165608
rect 580262 697176 580318 697232
rect 579618 683848 579674 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 579986 630808 580042 630864
rect 580170 617480 580226 617536
rect 580170 590960 580226 591016
rect 580170 577632 580226 577688
rect 580170 564304 580226 564360
rect 579894 537784 579950 537840
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 580170 471416 580226 471472
rect 580170 458088 580226 458144
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 579802 365064 579858 365120
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 579618 325216 579674 325272
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 578882 272176 578938 272232
rect 579986 258848 580042 258904
rect 580170 245520 580226 245576
rect 580354 524456 580410 524512
rect 580446 431568 580502 431624
rect 580262 233824 580318 233880
rect 579986 232328 580042 232384
rect 580170 219000 580226 219056
rect 579986 205672 580042 205728
rect 579710 192480 579766 192536
rect 580262 179152 580318 179208
rect 580170 165824 580226 165880
rect 580262 152632 580318 152688
rect 580262 139304 580318 139360
rect 580170 125976 580226 126032
rect 303618 43424 303674 43480
rect 309138 57160 309194 57216
rect 328458 58520 328514 58576
rect 332690 19896 332746 19952
rect 335358 40568 335414 40624
rect 338118 54440 338174 54496
rect 340970 53080 341026 53136
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580354 112784 580410 112840
rect 580262 19760 580318 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580257 697234 580323 697237
rect 583520 697234 584960 697324
rect 580257 697232 584960 697234
rect 580257 697176 580262 697232
rect 580318 697176 584960 697232
rect 580257 697174 584960 697176
rect 580257 697171 580323 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 579613 683906 579679 683909
rect 583520 683906 584960 683996
rect 579613 683904 584960 683906
rect 579613 683848 579618 683904
rect 579674 683848 584960 683904
rect 579613 683846 584960 683848
rect 579613 683843 579679 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 579889 537842 579955 537845
rect 583520 537842 584960 537932
rect 579889 537840 584960 537842
rect 579889 537784 579894 537840
rect 579950 537784 584960 537840
rect 579889 537782 584960 537784
rect 579889 537779 579955 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580349 524514 580415 524517
rect 583520 524514 584960 524604
rect 580349 524512 584960 524514
rect 580349 524456 580354 524512
rect 580410 524456 584960 524512
rect 580349 524454 584960 524456
rect 580349 524451 580415 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 2773 475690 2839 475693
rect -960 475688 2839 475690
rect -960 475632 2778 475688
rect 2834 475632 2839 475688
rect -960 475630 2839 475632
rect -960 475540 480 475630
rect 2773 475627 2839 475630
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3233 462634 3299 462637
rect -960 462632 3299 462634
rect -960 462576 3238 462632
rect 3294 462576 3299 462632
rect -960 462574 3299 462576
rect -960 462484 480 462574
rect 3233 462571 3299 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580441 431626 580507 431629
rect 583520 431626 584960 431716
rect 580441 431624 584960 431626
rect 580441 431568 580446 431624
rect 580502 431568 584960 431624
rect 580441 431566 584960 431568
rect 580441 431563 580507 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3601 371378 3667 371381
rect -960 371376 3667 371378
rect -960 371320 3606 371376
rect 3662 371320 3667 371376
rect -960 371318 3667 371320
rect -960 371228 480 371318
rect 3601 371315 3667 371318
rect 579797 365122 579863 365125
rect 583520 365122 584960 365212
rect 579797 365120 584960 365122
rect 579797 365064 579802 365120
rect 579858 365064 584960 365120
rect 579797 365062 584960 365064
rect 579797 365059 579863 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3509 358458 3575 358461
rect -960 358456 3575 358458
rect -960 358400 3514 358456
rect 3570 358400 3575 358456
rect -960 358398 3575 358400
rect -960 358308 480 358398
rect 3509 358395 3575 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 579613 325274 579679 325277
rect 583520 325274 584960 325364
rect 579613 325272 584960 325274
rect 579613 325216 579618 325272
rect 579674 325216 584960 325272
rect 579613 325214 584960 325216
rect 579613 325211 579679 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3693 306234 3759 306237
rect -960 306232 3759 306234
rect -960 306176 3698 306232
rect 3754 306176 3759 306232
rect -960 306174 3759 306176
rect -960 306084 480 306174
rect 3693 306171 3759 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3325 293178 3391 293181
rect -960 293176 3391 293178
rect -960 293120 3330 293176
rect 3386 293120 3391 293176
rect -960 293118 3391 293120
rect -960 293028 480 293118
rect 3325 293115 3391 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 578877 272234 578943 272237
rect 583520 272234 584960 272324
rect 578877 272232 584960 272234
rect 578877 272176 578882 272232
rect 578938 272176 584960 272232
rect 578877 272174 584960 272176
rect 578877 272171 578943 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3417 267202 3483 267205
rect -960 267200 3483 267202
rect -960 267144 3422 267200
rect 3478 267144 3483 267200
rect -960 267142 3483 267144
rect -960 267052 480 267142
rect 3417 267139 3483 267142
rect 579981 258906 580047 258909
rect 583520 258906 584960 258996
rect 579981 258904 584960 258906
rect 579981 258848 579986 258904
rect 580042 258848 584960 258904
rect 579981 258846 584960 258848
rect 579981 258843 580047 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 68318 252860 68324 252924
rect 68388 252922 68394 252924
rect 119153 252922 119219 252925
rect 68388 252920 119219 252922
rect 68388 252864 119158 252920
rect 119214 252864 119219 252920
rect 68388 252862 119219 252864
rect 68388 252860 68394 252862
rect 119153 252859 119219 252862
rect 68686 252724 68692 252788
rect 68756 252786 68762 252788
rect 123569 252786 123635 252789
rect 68756 252784 123635 252786
rect 68756 252728 123574 252784
rect 123630 252728 123635 252784
rect 68756 252726 123635 252728
rect 68756 252724 68762 252726
rect 123569 252723 123635 252726
rect 68502 252588 68508 252652
rect 68572 252650 68578 252652
rect 123753 252650 123819 252653
rect 68572 252648 123819 252650
rect 68572 252592 123758 252648
rect 123814 252592 123819 252648
rect 68572 252590 123819 252592
rect 68572 252588 68578 252590
rect 123753 252587 123819 252590
rect 106089 251970 106155 251973
rect 120022 251970 120028 251972
rect 106089 251968 120028 251970
rect 106089 251912 106094 251968
rect 106150 251912 120028 251968
rect 106089 251910 120028 251912
rect 106089 251907 106155 251910
rect 120022 251908 120028 251910
rect 120092 251908 120098 251972
rect 69054 251772 69060 251836
rect 69124 251834 69130 251836
rect 71957 251834 72023 251837
rect 73061 251834 73127 251837
rect 119889 251834 119955 251837
rect 69124 251832 119955 251834
rect 69124 251776 71962 251832
rect 72018 251776 73066 251832
rect 73122 251776 119894 251832
rect 119950 251776 119955 251832
rect 69124 251774 119955 251776
rect 69124 251772 69130 251774
rect 71957 251771 72023 251774
rect 73061 251771 73127 251774
rect 119889 251771 119955 251774
rect 94681 251698 94747 251701
rect 119245 251698 119311 251701
rect 94681 251696 119311 251698
rect 94681 251640 94686 251696
rect 94742 251640 119250 251696
rect 119306 251640 119311 251696
rect 94681 251638 119311 251640
rect 94681 251635 94747 251638
rect 119245 251635 119311 251638
rect 65977 251562 66043 251565
rect 84193 251562 84259 251565
rect 119838 251562 119844 251564
rect 65977 251560 119844 251562
rect 65977 251504 65982 251560
rect 66038 251504 84198 251560
rect 84254 251504 119844 251560
rect 65977 251502 119844 251504
rect 65977 251499 66043 251502
rect 84193 251499 84259 251502
rect 119838 251500 119844 251502
rect 119908 251500 119914 251564
rect 64689 251426 64755 251429
rect 84837 251426 84903 251429
rect 118693 251426 118759 251429
rect 64689 251424 118759 251426
rect 64689 251368 64694 251424
rect 64750 251368 84842 251424
rect 84898 251368 118698 251424
rect 118754 251368 118759 251424
rect 64689 251366 118759 251368
rect 64689 251363 64755 251366
rect 84837 251363 84903 251366
rect 118693 251363 118759 251366
rect 116393 251290 116459 251293
rect 131113 251290 131179 251293
rect 116393 251288 131179 251290
rect 116393 251232 116398 251288
rect 116454 251232 131118 251288
rect 131174 251232 131179 251288
rect 116393 251230 131179 251232
rect 116393 251227 116459 251230
rect 131113 251227 131179 251230
rect 103421 251154 103487 251157
rect 103421 251152 113190 251154
rect 103421 251096 103426 251152
rect 103482 251096 113190 251152
rect 103421 251094 113190 251096
rect 103421 251091 103487 251094
rect 113130 250610 113190 251094
rect 152457 250610 152523 250613
rect 113130 250608 152523 250610
rect 113130 250552 152462 250608
rect 152518 250552 152523 250608
rect 113130 250550 152523 250552
rect 152457 250547 152523 250550
rect 95141 250474 95207 250477
rect 178033 250474 178099 250477
rect 95141 250472 178099 250474
rect 95141 250416 95146 250472
rect 95202 250416 178038 250472
rect 178094 250416 178099 250472
rect 95141 250414 178099 250416
rect 95141 250411 95207 250414
rect 178033 250411 178099 250414
rect 88701 250202 88767 250205
rect 119470 250202 119476 250204
rect 88701 250200 119476 250202
rect 88701 250144 88706 250200
rect 88762 250144 119476 250200
rect 88701 250142 119476 250144
rect 88701 250139 88767 250142
rect 119470 250140 119476 250142
rect 119540 250140 119546 250204
rect 82261 250066 82327 250069
rect 119654 250066 119660 250068
rect 82261 250064 119660 250066
rect 82261 250008 82266 250064
rect 82322 250008 119660 250064
rect 82261 250006 119660 250008
rect 82261 250003 82327 250006
rect 119654 250004 119660 250006
rect 119724 250004 119730 250068
rect 78397 249930 78463 249933
rect 119337 249930 119403 249933
rect 78397 249928 119403 249930
rect 78397 249872 78402 249928
rect 78458 249872 119342 249928
rect 119398 249872 119403 249928
rect 78397 249870 119403 249872
rect 78397 249867 78463 249870
rect 119337 249867 119403 249870
rect 68737 249794 68803 249797
rect 112161 249794 112227 249797
rect 182173 249794 182239 249797
rect 182817 249794 182883 249797
rect 68737 249792 70380 249794
rect 68737 249736 68742 249792
rect 68798 249736 70380 249792
rect 68737 249734 70380 249736
rect 112161 249792 182883 249794
rect 112161 249736 112166 249792
rect 112222 249736 182178 249792
rect 182234 249736 182822 249792
rect 182878 249736 182883 249792
rect 112161 249734 182883 249736
rect 68737 249731 68803 249734
rect 112161 249731 112227 249734
rect 182173 249731 182239 249734
rect 182817 249731 182883 249734
rect 122373 248978 122439 248981
rect 119692 248976 122439 248978
rect 119692 248920 122378 248976
rect 122434 248920 122439 248976
rect 119692 248918 122439 248920
rect 122373 248915 122439 248918
rect 68829 248300 68895 248301
rect 68829 248298 68876 248300
rect 68748 248296 68876 248298
rect 68940 248298 68946 248300
rect 121453 248298 121519 248301
rect 68748 248240 68834 248296
rect 68748 248238 68876 248240
rect 68829 248236 68876 248238
rect 68940 248238 70380 248298
rect 119692 248296 121519 248298
rect 119692 248240 121458 248296
rect 121514 248240 121519 248296
rect 119692 248238 121519 248240
rect 68940 248236 68946 248238
rect 68829 248235 68895 248236
rect 121453 248235 121519 248238
rect 119838 247964 119844 248028
rect 119908 248026 119914 248028
rect 187049 248026 187115 248029
rect 119908 248024 187115 248026
rect 119908 247968 187054 248024
rect 187110 247968 187115 248024
rect 119908 247966 187115 247968
rect 119908 247964 119914 247966
rect 187049 247963 187115 247966
rect 67633 247754 67699 247757
rect 68553 247754 68619 247757
rect 67633 247752 70380 247754
rect 67633 247696 67638 247752
rect 67694 247696 68558 247752
rect 68614 247696 70380 247752
rect 67633 247694 70380 247696
rect 67633 247691 67699 247694
rect 68553 247691 68619 247694
rect 120022 247556 120028 247620
rect 120092 247618 120098 247620
rect 133137 247618 133203 247621
rect 133781 247618 133847 247621
rect 120092 247616 133847 247618
rect 120092 247560 133142 247616
rect 133198 247560 133786 247616
rect 133842 247560 133847 247616
rect 120092 247558 133847 247560
rect 120092 247556 120098 247558
rect 133137 247555 133203 247558
rect 133781 247555 133847 247558
rect 121453 246938 121519 246941
rect 119692 246936 121519 246938
rect 119692 246880 121458 246936
rect 121514 246880 121519 246936
rect 119692 246878 121519 246880
rect 121453 246875 121519 246878
rect 69105 246258 69171 246261
rect 69105 246256 70380 246258
rect 69105 246200 69110 246256
rect 69166 246200 70380 246256
rect 69105 246198 70380 246200
rect 69105 246195 69171 246198
rect 119662 245850 119722 246228
rect 121862 246196 121868 246260
rect 121932 246258 121938 246260
rect 122005 246258 122071 246261
rect 121932 246256 122071 246258
rect 121932 246200 122010 246256
rect 122066 246200 122071 246256
rect 121932 246198 122071 246200
rect 121932 246196 121938 246198
rect 122005 246195 122071 246198
rect 122649 245850 122715 245853
rect 119662 245848 122715 245850
rect 119662 245792 122654 245848
rect 122710 245792 122715 245848
rect 119662 245790 122715 245792
rect 122649 245787 122715 245790
rect 67541 245578 67607 245581
rect 68277 245578 68343 245581
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 67541 245576 70380 245578
rect 67541 245520 67546 245576
rect 67602 245520 68282 245576
rect 68338 245520 70380 245576
rect 67541 245518 70380 245520
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 67541 245515 67607 245518
rect 68277 245515 68343 245518
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 121637 244898 121703 244901
rect 119692 244896 121703 244898
rect 119692 244840 121642 244896
rect 121698 244840 121703 244896
rect 119692 244838 121703 244840
rect 121637 244835 121703 244838
rect 67633 244354 67699 244357
rect 121453 244354 121519 244357
rect 67633 244352 70380 244354
rect 67633 244296 67638 244352
rect 67694 244296 70380 244352
rect 67633 244294 70380 244296
rect 119692 244352 121519 244354
rect 119692 244296 121458 244352
rect 121514 244296 121519 244352
rect 119692 244294 121519 244296
rect 67633 244291 67699 244294
rect 121453 244291 121519 244294
rect 68645 243674 68711 243677
rect 68645 243672 68754 243674
rect 68645 243616 68650 243672
rect 68706 243616 68754 243672
rect 68645 243611 68754 243616
rect 68694 243402 68754 243611
rect 69473 243538 69539 243541
rect 69473 243536 70380 243538
rect 69473 243480 69478 243536
rect 69534 243480 70380 243536
rect 69473 243478 70380 243480
rect 69473 243475 69539 243478
rect 68694 243342 70410 243402
rect 70350 242964 70410 243342
rect 122281 242996 122347 242997
rect 122230 242994 122236 242996
rect 119692 242934 122236 242994
rect 122300 242994 122347 242996
rect 122300 242992 122392 242994
rect 122342 242936 122392 242992
rect 122230 242932 122236 242934
rect 122300 242934 122392 242936
rect 122300 242932 122347 242934
rect 122281 242931 122347 242932
rect 121453 242178 121519 242181
rect 119692 242176 121519 242178
rect 119692 242120 121458 242176
rect 121514 242120 121519 242176
rect 119692 242118 121519 242120
rect 121453 242115 121519 242118
rect 67214 241572 67220 241636
rect 67284 241634 67290 241636
rect 67449 241634 67515 241637
rect 121545 241634 121611 241637
rect 67284 241632 70380 241634
rect 67284 241576 67454 241632
rect 67510 241576 70380 241632
rect 67284 241574 70380 241576
rect 119692 241632 121611 241634
rect 119692 241576 121550 241632
rect 121606 241576 121611 241632
rect 119692 241574 121611 241576
rect 67284 241572 67290 241574
rect 67449 241571 67515 241574
rect 121545 241571 121611 241574
rect -960 241090 480 241180
rect 3049 241090 3115 241093
rect -960 241088 3115 241090
rect -960 241032 3054 241088
rect 3110 241032 3115 241088
rect -960 241030 3115 241032
rect -960 240940 480 241030
rect 3049 241027 3115 241030
rect 68369 240954 68435 240957
rect 68369 240952 70380 240954
rect 68369 240896 68374 240952
rect 68430 240896 70380 240952
rect 68369 240894 70380 240896
rect 68369 240891 68435 240894
rect 120206 240274 120212 240276
rect 119692 240214 120212 240274
rect 120206 240212 120212 240214
rect 120276 240274 120282 240276
rect 230422 240274 230428 240276
rect 120276 240214 230428 240274
rect 120276 240212 120282 240214
rect 230422 240212 230428 240214
rect 230492 240212 230498 240276
rect 68318 239532 68324 239596
rect 68388 239594 68394 239596
rect 121821 239594 121887 239597
rect 68388 239534 70380 239594
rect 119692 239592 121887 239594
rect 119692 239536 121826 239592
rect 121882 239536 121887 239592
rect 119692 239534 121887 239536
rect 68388 239532 68394 239534
rect 121821 239531 121887 239534
rect 68502 238852 68508 238916
rect 68572 238914 68578 238916
rect 68572 238854 70380 238914
rect 68572 238852 68578 238854
rect 121453 238098 121519 238101
rect 119692 238096 121519 238098
rect 119692 238040 121458 238096
rect 121514 238040 121519 238096
rect 119692 238038 121519 238040
rect 121453 238035 121519 238038
rect 68829 237554 68895 237557
rect 68829 237552 70380 237554
rect 68829 237496 68834 237552
rect 68890 237496 70380 237552
rect 68829 237494 70380 237496
rect 68829 237491 68895 237494
rect 121821 237418 121887 237421
rect 119692 237416 121887 237418
rect 119692 237360 121826 237416
rect 121882 237360 121887 237416
rect 119692 237358 121887 237360
rect 121821 237355 121887 237358
rect 68369 236874 68435 236877
rect 68369 236872 70380 236874
rect 68369 236816 68374 236872
rect 68430 236816 70380 236872
rect 68369 236814 70380 236816
rect 68369 236811 68435 236814
rect 69381 236194 69447 236197
rect 69381 236192 70380 236194
rect 69381 236136 69386 236192
rect 69442 236136 70380 236192
rect 69381 236134 70380 236136
rect 69381 236131 69447 236134
rect 122741 236058 122807 236061
rect 119692 236056 122807 236058
rect 119692 236000 122746 236056
rect 122802 236000 122807 236056
rect 119692 235998 122807 236000
rect 122741 235995 122807 235998
rect 122281 235378 122347 235381
rect 119692 235376 122347 235378
rect 119692 235320 122286 235376
rect 122342 235320 122347 235376
rect 119692 235318 122347 235320
rect 122281 235315 122347 235318
rect 69289 234834 69355 234837
rect 69289 234832 70380 234834
rect 69289 234776 69294 234832
rect 69350 234776 70380 234832
rect 69289 234774 70380 234776
rect 69289 234771 69355 234774
rect 122465 234698 122531 234701
rect 119692 234696 122531 234698
rect 119692 234640 122470 234696
rect 122526 234640 122531 234696
rect 119692 234638 122531 234640
rect 122465 234635 122531 234638
rect 69013 234154 69079 234157
rect 69013 234152 70380 234154
rect 69013 234096 69018 234152
rect 69074 234096 70380 234152
rect 69013 234094 70380 234096
rect 69013 234091 69079 234094
rect 169518 233820 169524 233884
rect 169588 233882 169594 233884
rect 580257 233882 580323 233885
rect 169588 233880 580323 233882
rect 169588 233824 580262 233880
rect 580318 233824 580323 233880
rect 169588 233822 580323 233824
rect 169588 233820 169594 233822
rect 580257 233819 580323 233822
rect 122465 233338 122531 233341
rect 119692 233336 122531 233338
rect 119692 233280 122470 233336
rect 122526 233280 122531 233336
rect 119692 233278 122531 233280
rect 122465 233275 122531 233278
rect 183553 233202 183619 233205
rect 184197 233202 184263 233205
rect 122790 233200 184263 233202
rect 122790 233144 183558 233200
rect 183614 233144 184202 233200
rect 184258 233144 184263 233200
rect 122790 233142 184263 233144
rect 119838 233004 119844 233068
rect 119908 233066 119914 233068
rect 122790 233066 122850 233142
rect 183553 233139 183619 233142
rect 184197 233139 184263 233142
rect 119908 233006 122850 233066
rect 119908 233004 119914 233006
rect 121729 232794 121795 232797
rect 119692 232792 121795 232794
rect 119692 232736 121734 232792
rect 121790 232736 121795 232792
rect 119692 232734 121795 232736
rect 121729 232731 121795 232734
rect 68737 232660 68803 232661
rect 68686 232658 68692 232660
rect 68610 232598 68692 232658
rect 68756 232658 68803 232660
rect 68756 232656 70380 232658
rect 68798 232600 70380 232656
rect 68686 232596 68692 232598
rect 68756 232598 70380 232600
rect 68756 232596 68803 232598
rect 68737 232595 68803 232596
rect 119470 232460 119476 232524
rect 119540 232522 119546 232524
rect 140773 232522 140839 232525
rect 119540 232520 140839 232522
rect 119540 232464 140778 232520
rect 140834 232464 140839 232520
rect 119540 232462 140839 232464
rect 119540 232460 119546 232462
rect 140773 232459 140839 232462
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect 68369 232114 68435 232117
rect 68369 232112 70380 232114
rect 68369 232056 68374 232112
rect 68430 232056 70380 232112
rect 68369 232054 70380 232056
rect 68369 232051 68435 232054
rect 119294 231029 119354 231268
rect 119294 231024 119403 231029
rect 119294 230968 119342 231024
rect 119398 230968 119403 231024
rect 119294 230966 119403 230968
rect 119337 230963 119403 230966
rect 121453 230754 121519 230757
rect 119692 230752 121519 230754
rect 119692 230696 121458 230752
rect 121514 230696 121519 230752
rect 119692 230694 121519 230696
rect 121453 230691 121519 230694
rect 67633 230618 67699 230621
rect 67633 230616 70380 230618
rect 67633 230560 67638 230616
rect 67694 230560 70380 230616
rect 67633 230558 70380 230560
rect 67633 230555 67699 230558
rect 169702 230556 169708 230620
rect 169772 230618 169778 230620
rect 171225 230618 171291 230621
rect 169772 230616 171291 230618
rect 169772 230560 171230 230616
rect 171286 230560 171291 230616
rect 169772 230558 171291 230560
rect 169772 230556 169778 230558
rect 171225 230555 171291 230558
rect 68645 230074 68711 230077
rect 68645 230072 70380 230074
rect 68645 230016 68650 230072
rect 68706 230016 70380 230072
rect 68645 230014 70380 230016
rect 68645 230011 68711 230014
rect 67725 229394 67791 229397
rect 67725 229392 70380 229394
rect 67725 229336 67730 229392
rect 67786 229336 70380 229392
rect 67725 229334 70380 229336
rect 67725 229331 67791 229334
rect 119654 229196 119660 229260
rect 119724 229258 119730 229260
rect 121453 229258 121519 229261
rect 119724 229256 121519 229258
rect 119724 229200 121458 229256
rect 121514 229200 121519 229256
rect 119724 229198 121519 229200
rect 119724 229196 119730 229198
rect 121453 229195 121519 229198
rect 166993 229258 167059 229261
rect 166993 229256 170292 229258
rect 166993 229200 166998 229256
rect 167054 229200 170292 229256
rect 166993 229198 170292 229200
rect 166993 229195 167059 229198
rect 229326 229062 229754 229122
rect 229326 228986 229386 229062
rect 119294 228926 229386 228986
rect 229694 228986 229754 229062
rect 229829 228986 229895 228989
rect 229694 228984 229895 228986
rect 229694 228928 229834 228984
rect 229890 228928 229895 228984
rect 229694 228926 229895 228928
rect 119294 228580 119354 228926
rect 229829 228923 229895 228926
rect 229277 228850 229343 228853
rect 122790 228848 229343 228850
rect 122790 228792 229282 228848
rect 229338 228792 229343 228848
rect 122790 228790 229343 228792
rect 119286 228516 119292 228580
rect 119356 228516 119362 228580
rect 122790 228442 122850 228790
rect 229277 228787 229343 228790
rect 229461 228850 229527 228853
rect 229461 228848 229570 228850
rect 229461 228792 229466 228848
rect 229522 228792 229570 228848
rect 229461 228787 229570 228792
rect 229510 228548 229570 228787
rect 119662 228382 122850 228442
rect -960 227884 480 228124
rect 68461 228034 68527 228037
rect 68461 228032 70380 228034
rect 68461 227976 68466 228032
rect 68522 227976 70380 228032
rect 68461 227974 70380 227976
rect 68461 227971 68527 227974
rect 119662 227898 119722 228382
rect 120022 227898 120028 227900
rect 119662 227868 120028 227898
rect 119692 227838 120028 227868
rect 120022 227836 120028 227838
rect 120092 227836 120098 227900
rect 167085 227898 167151 227901
rect 167085 227896 170292 227898
rect 167085 227840 167090 227896
rect 167146 227840 170292 227896
rect 167085 227838 170292 227840
rect 167085 227835 167151 227838
rect 229277 227762 229343 227765
rect 231894 227762 231900 227764
rect 229277 227760 231900 227762
rect 229277 227704 229282 227760
rect 229338 227704 231900 227760
rect 229277 227702 231900 227704
rect 229277 227699 229343 227702
rect 231894 227700 231900 227702
rect 231964 227700 231970 227764
rect 68921 227354 68987 227357
rect 68921 227352 70380 227354
rect 68921 227296 68926 227352
rect 68982 227296 70380 227352
rect 68921 227294 70380 227296
rect 68921 227291 68987 227294
rect 167545 227218 167611 227221
rect 230289 227218 230355 227221
rect 167545 227216 170292 227218
rect 167545 227160 167550 227216
rect 167606 227160 170292 227216
rect 229724 227216 230355 227218
rect 229724 227188 230294 227216
rect 167545 227158 170292 227160
rect 229694 227160 230294 227188
rect 230350 227160 230355 227216
rect 229694 227158 230355 227160
rect 167545 227155 167611 227158
rect 229694 226677 229754 227158
rect 230289 227155 230355 227158
rect 229645 226672 229754 226677
rect 229645 226616 229650 226672
rect 229706 226616 229754 226672
rect 229645 226614 229754 226616
rect 229645 226611 229711 226614
rect 119662 226402 119722 226508
rect 120574 226402 120580 226404
rect 119662 226342 120580 226402
rect 120574 226340 120580 226342
rect 120644 226340 120650 226404
rect 67817 225858 67883 225861
rect 68185 225858 68251 225861
rect 122465 225858 122531 225861
rect 67817 225856 70380 225858
rect 67817 225800 67822 225856
rect 67878 225800 68190 225856
rect 68246 225800 70380 225856
rect 67817 225798 70380 225800
rect 119692 225856 122531 225858
rect 119692 225800 122470 225856
rect 122526 225800 122531 225856
rect 119692 225798 122531 225800
rect 67817 225795 67883 225798
rect 68185 225795 68251 225798
rect 122465 225795 122531 225798
rect 167085 225858 167151 225861
rect 230197 225858 230263 225861
rect 167085 225856 170292 225858
rect 167085 225800 167090 225856
rect 167146 225800 170292 225856
rect 167085 225798 170292 225800
rect 229724 225856 230263 225858
rect 229724 225800 230202 225856
rect 230258 225800 230263 225856
rect 229724 225798 230263 225800
rect 167085 225795 167151 225798
rect 230197 225795 230263 225798
rect 68737 225314 68803 225317
rect 69013 225314 69079 225317
rect 68737 225312 70380 225314
rect 68737 225256 68742 225312
rect 68798 225256 69018 225312
rect 69074 225256 70380 225312
rect 68737 225254 70380 225256
rect 68737 225251 68803 225254
rect 69013 225251 69079 225254
rect 232681 225178 232747 225181
rect 229724 225176 232747 225178
rect 229724 225120 232686 225176
rect 232742 225120 232747 225176
rect 229724 225118 232747 225120
rect 232681 225115 232747 225118
rect 121453 224634 121519 224637
rect 119692 224632 121519 224634
rect 119692 224576 121458 224632
rect 121514 224576 121519 224632
rect 119692 224574 121519 224576
rect 121453 224571 121519 224574
rect 167085 224498 167151 224501
rect 167085 224496 170292 224498
rect 167085 224440 167090 224496
rect 167146 224440 170292 224496
rect 167085 224438 170292 224440
rect 167085 224435 167151 224438
rect 66897 223818 66963 223821
rect 122189 223818 122255 223821
rect 231301 223818 231367 223821
rect 66897 223816 70380 223818
rect 66897 223760 66902 223816
rect 66958 223760 70380 223816
rect 66897 223758 70380 223760
rect 119692 223816 122255 223818
rect 119692 223760 122194 223816
rect 122250 223760 122255 223816
rect 119692 223758 122255 223760
rect 229724 223816 231367 223818
rect 229724 223760 231306 223816
rect 231362 223760 231367 223816
rect 229724 223758 231367 223760
rect 66897 223755 66963 223758
rect 122189 223755 122255 223758
rect 231301 223755 231367 223758
rect 68645 223138 68711 223141
rect 167085 223138 167151 223141
rect 68645 223136 70380 223138
rect 68645 223080 68650 223136
rect 68706 223080 70380 223136
rect 68645 223078 70380 223080
rect 167085 223136 170292 223138
rect 167085 223080 167090 223136
rect 167146 223080 170292 223136
rect 167085 223078 170292 223080
rect 68645 223075 68711 223078
rect 167085 223075 167151 223078
rect 121545 222594 121611 222597
rect 121913 222594 121979 222597
rect 119692 222592 121979 222594
rect 119692 222536 121550 222592
rect 121606 222536 121918 222592
rect 121974 222536 121979 222592
rect 119692 222534 121979 222536
rect 121545 222531 121611 222534
rect 121913 222531 121979 222534
rect 167821 222458 167887 222461
rect 230933 222458 230999 222461
rect 167821 222456 170292 222458
rect 167821 222400 167826 222456
rect 167882 222400 170292 222456
rect 167821 222398 170292 222400
rect 229724 222456 230999 222458
rect 229724 222400 230938 222456
rect 230994 222400 230999 222456
rect 229724 222398 230999 222400
rect 167821 222395 167887 222398
rect 230933 222395 230999 222398
rect 121453 221914 121519 221917
rect 119692 221912 121519 221914
rect 119692 221884 121458 221912
rect 119662 221856 121458 221884
rect 121514 221856 121519 221912
rect 119662 221854 121519 221856
rect 69473 221778 69539 221781
rect 69473 221776 70380 221778
rect 69473 221720 69478 221776
rect 69534 221720 70380 221776
rect 69473 221718 70380 221720
rect 69473 221715 69539 221718
rect 119286 221172 119292 221236
rect 119356 221234 119362 221236
rect 119662 221234 119722 221854
rect 121453 221851 121519 221854
rect 119356 221174 119722 221234
rect 119356 221172 119362 221174
rect 68001 221098 68067 221101
rect 167453 221098 167519 221101
rect 230105 221098 230171 221101
rect 68001 221096 70380 221098
rect 68001 221040 68006 221096
rect 68062 221040 70380 221096
rect 68001 221038 70380 221040
rect 167453 221096 170292 221098
rect 167453 221040 167458 221096
rect 167514 221040 170292 221096
rect 167453 221038 170292 221040
rect 229724 221096 230171 221098
rect 229724 221040 230110 221096
rect 230166 221040 230171 221096
rect 229724 221038 230171 221040
rect 68001 221035 68067 221038
rect 167453 221035 167519 221038
rect 230105 221035 230171 221038
rect 68921 220418 68987 220421
rect 120441 220418 120507 220421
rect 231393 220418 231459 220421
rect 68921 220416 70380 220418
rect 68921 220360 68926 220416
rect 68982 220360 70380 220416
rect 68921 220358 70380 220360
rect 119692 220416 120507 220418
rect 119692 220360 120446 220416
rect 120502 220360 120507 220416
rect 119692 220358 120507 220360
rect 229724 220416 231459 220418
rect 229724 220360 231398 220416
rect 231454 220360 231459 220416
rect 229724 220358 231459 220360
rect 68921 220355 68987 220358
rect 120441 220355 120507 220358
rect 231393 220355 231459 220358
rect 120165 219874 120231 219877
rect 119692 219872 120231 219874
rect 119692 219844 120170 219872
rect 119662 219816 120170 219844
rect 120226 219816 120231 219872
rect 119662 219814 120231 219816
rect 119337 219602 119403 219605
rect 119662 219602 119722 219814
rect 120165 219811 120231 219814
rect 167729 219738 167795 219741
rect 167729 219736 170292 219738
rect 167729 219680 167734 219736
rect 167790 219680 170292 219736
rect 167729 219678 170292 219680
rect 167729 219675 167795 219678
rect 119337 219600 119722 219602
rect 119337 219544 119342 219600
rect 119398 219544 119722 219600
rect 119337 219542 119722 219544
rect 119337 219539 119403 219542
rect 68185 219058 68251 219061
rect 167085 219058 167151 219061
rect 230013 219058 230079 219061
rect 68185 219056 70380 219058
rect 68185 219000 68190 219056
rect 68246 219000 70380 219056
rect 167085 219056 170292 219058
rect 68185 218998 70380 219000
rect 68185 218995 68251 218998
rect 119478 218517 119538 219028
rect 167085 219000 167090 219056
rect 167146 219000 170292 219056
rect 167085 218998 170292 219000
rect 229724 219056 230079 219058
rect 229724 219000 230018 219056
rect 230074 219000 230079 219056
rect 229724 218998 230079 219000
rect 167085 218995 167151 218998
rect 230013 218995 230079 218998
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect 119478 218512 119587 218517
rect 119478 218456 119526 218512
rect 119582 218456 119587 218512
rect 119478 218454 119587 218456
rect 119521 218451 119587 218454
rect 68461 218378 68527 218381
rect 68461 218376 70380 218378
rect 68461 218320 68466 218376
rect 68522 218320 70380 218376
rect 68461 218318 70380 218320
rect 68461 218315 68527 218318
rect 230422 217970 230428 217972
rect 229694 217910 230428 217970
rect 120165 217698 120231 217701
rect 119692 217696 120231 217698
rect 119692 217640 120170 217696
rect 120226 217640 120231 217696
rect 119692 217638 120231 217640
rect 120165 217635 120231 217638
rect 167085 217698 167151 217701
rect 167494 217698 167500 217700
rect 167085 217696 167500 217698
rect 167085 217640 167090 217696
rect 167146 217640 167500 217696
rect 167085 217638 167500 217640
rect 167085 217635 167151 217638
rect 167494 217636 167500 217638
rect 167564 217698 167570 217700
rect 167564 217638 170292 217698
rect 229694 217668 229754 217910
rect 230422 217908 230428 217910
rect 230492 217970 230498 217972
rect 232681 217970 232747 217973
rect 230492 217968 232747 217970
rect 230492 217912 232686 217968
rect 232742 217912 232747 217968
rect 230492 217910 232747 217912
rect 230492 217908 230498 217910
rect 232681 217907 232747 217910
rect 167564 217636 167570 217638
rect 68369 217018 68435 217021
rect 122005 217018 122071 217021
rect 231209 217018 231275 217021
rect 68369 217016 70380 217018
rect 68369 216960 68374 217016
rect 68430 216960 70380 217016
rect 68369 216958 70380 216960
rect 119692 217016 122071 217018
rect 119692 216960 122010 217016
rect 122066 216960 122071 217016
rect 119692 216958 122071 216960
rect 229724 217016 231275 217018
rect 229724 216960 231214 217016
rect 231270 216960 231275 217016
rect 229724 216958 231275 216960
rect 68369 216955 68435 216958
rect 122005 216955 122071 216958
rect 231209 216955 231275 216958
rect 67633 216338 67699 216341
rect 167085 216338 167151 216341
rect 67633 216336 70380 216338
rect 67633 216280 67638 216336
rect 67694 216280 70380 216336
rect 67633 216278 70380 216280
rect 167085 216336 170292 216338
rect 167085 216280 167090 216336
rect 167146 216280 170292 216336
rect 167085 216278 170292 216280
rect 67633 216275 67699 216278
rect 167085 216275 167151 216278
rect 121453 215794 121519 215797
rect 119692 215792 121519 215794
rect 119692 215736 121458 215792
rect 121514 215736 121519 215792
rect 119692 215734 121519 215736
rect 121453 215731 121519 215734
rect 231117 215658 231183 215661
rect 229724 215656 231183 215658
rect 229724 215600 231122 215656
rect 231178 215600 231183 215656
rect 229724 215598 231183 215600
rect 231117 215595 231183 215598
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 68369 214978 68435 214981
rect 121453 214978 121519 214981
rect 68369 214976 70380 214978
rect 68369 214920 68374 214976
rect 68430 214920 70380 214976
rect 68369 214918 70380 214920
rect 119692 214976 121519 214978
rect 119692 214920 121458 214976
rect 121514 214920 121519 214976
rect 119692 214918 121519 214920
rect 68369 214915 68435 214918
rect 121453 214915 121519 214918
rect 167177 214978 167243 214981
rect 167177 214976 170292 214978
rect 167177 214920 167182 214976
rect 167238 214920 170292 214976
rect 167177 214918 170292 214920
rect 167177 214915 167243 214918
rect 67633 214434 67699 214437
rect 68185 214434 68251 214437
rect 67633 214432 70380 214434
rect 67633 214376 67638 214432
rect 67694 214376 68190 214432
rect 68246 214376 70380 214432
rect 67633 214374 70380 214376
rect 67633 214371 67699 214374
rect 68185 214371 68251 214374
rect 167085 214298 167151 214301
rect 230749 214298 230815 214301
rect 167085 214296 170292 214298
rect 167085 214240 167090 214296
rect 167146 214240 170292 214296
rect 167085 214238 170292 214240
rect 229724 214296 230815 214298
rect 229724 214240 230754 214296
rect 230810 214240 230815 214296
rect 229724 214238 230815 214240
rect 167085 214235 167151 214238
rect 230749 214235 230815 214238
rect 67909 213618 67975 213621
rect 121913 213618 121979 213621
rect 67909 213616 70380 213618
rect 67909 213560 67914 213616
rect 67970 213560 70380 213616
rect 67909 213558 70380 213560
rect 119692 213616 121979 213618
rect 119692 213560 121918 213616
rect 121974 213560 121979 213616
rect 119692 213558 121979 213560
rect 67909 213555 67975 213558
rect 121913 213555 121979 213558
rect 121729 213074 121795 213077
rect 122046 213074 122052 213076
rect 119692 213072 122052 213074
rect 119692 213016 121734 213072
rect 121790 213016 122052 213072
rect 119692 213014 122052 213016
rect 121729 213011 121795 213014
rect 122046 213012 122052 213014
rect 122116 213012 122122 213076
rect 167637 212938 167703 212941
rect 230565 212938 230631 212941
rect 167637 212936 170292 212938
rect 167637 212880 167642 212936
rect 167698 212880 170292 212936
rect 167637 212878 170292 212880
rect 229724 212936 230631 212938
rect 229724 212880 230570 212936
rect 230626 212880 230631 212936
rect 229724 212878 230631 212880
rect 167637 212875 167703 212878
rect 230565 212875 230631 212878
rect 229553 212530 229619 212533
rect 229510 212528 229619 212530
rect 229510 212472 229558 212528
rect 229614 212472 229619 212528
rect 229510 212467 229619 212472
rect 121453 212258 121519 212261
rect 119692 212256 121519 212258
rect 69657 211986 69723 211989
rect 70350 211986 70410 212228
rect 119692 212200 121458 212256
rect 121514 212200 121519 212256
rect 229510 212258 229570 212467
rect 230565 212258 230631 212261
rect 229510 212256 230631 212258
rect 229510 212228 230570 212256
rect 119692 212198 121519 212200
rect 229540 212200 230570 212228
rect 230626 212200 230631 212256
rect 229540 212198 230631 212200
rect 121453 212195 121519 212198
rect 230565 212195 230631 212198
rect 69657 211984 70410 211986
rect 69657 211928 69662 211984
rect 69718 211928 70410 211984
rect 69657 211926 70410 211928
rect 69657 211923 69723 211926
rect 69381 211578 69447 211581
rect 167085 211578 167151 211581
rect 167361 211578 167427 211581
rect 69381 211576 70380 211578
rect 69381 211520 69386 211576
rect 69442 211520 70380 211576
rect 69381 211518 70380 211520
rect 167085 211576 170292 211578
rect 167085 211520 167090 211576
rect 167146 211520 167366 211576
rect 167422 211520 170292 211576
rect 167085 211518 170292 211520
rect 69381 211515 69447 211518
rect 167085 211515 167151 211518
rect 167361 211515 167427 211518
rect 121545 211034 121611 211037
rect 119692 211032 121611 211034
rect 119692 211004 121550 211032
rect 119662 210976 121550 211004
rect 121606 210976 121611 211032
rect 119662 210974 121611 210976
rect 119286 210700 119292 210764
rect 119356 210762 119362 210764
rect 119662 210762 119722 210974
rect 121545 210971 121611 210974
rect 167085 210898 167151 210901
rect 167269 210898 167335 210901
rect 230473 210898 230539 210901
rect 167085 210896 170292 210898
rect 167085 210840 167090 210896
rect 167146 210840 167274 210896
rect 167330 210840 170292 210896
rect 167085 210838 170292 210840
rect 229724 210896 230539 210898
rect 229724 210840 230478 210896
rect 230534 210840 230539 210896
rect 229724 210838 230539 210840
rect 167085 210835 167151 210838
rect 167269 210835 167335 210838
rect 230473 210835 230539 210838
rect 119356 210702 119722 210762
rect 119356 210700 119362 210702
rect 65333 210218 65399 210221
rect 68686 210218 68692 210220
rect 65333 210216 68692 210218
rect 65333 210160 65338 210216
rect 65394 210160 68692 210216
rect 65333 210158 68692 210160
rect 65333 210155 65399 210158
rect 68686 210156 68692 210158
rect 68756 210218 68762 210220
rect 122414 210218 122420 210220
rect 68756 210158 70380 210218
rect 119692 210158 122420 210218
rect 68756 210156 68762 210158
rect 122414 210156 122420 210158
rect 122484 210156 122490 210220
rect 70710 209476 70716 209540
rect 70780 209476 70786 209540
rect 168189 209538 168255 209541
rect 230381 209538 230447 209541
rect 168189 209536 170292 209538
rect 168189 209480 168194 209536
rect 168250 209480 170292 209536
rect 168189 209478 170292 209480
rect 229724 209536 230447 209538
rect 229724 209480 230386 209536
rect 230442 209480 230447 209536
rect 229724 209478 230447 209480
rect 168189 209475 168255 209478
rect 230381 209475 230447 209478
rect 229277 209266 229343 209269
rect 229277 209264 229386 209266
rect 229277 209208 229282 209264
rect 229338 209208 229386 209264
rect 229277 209203 229386 209208
rect 122373 208858 122439 208861
rect 119692 208856 122439 208858
rect 119692 208800 122378 208856
rect 122434 208800 122439 208856
rect 229326 208828 229386 209203
rect 119692 208798 122439 208800
rect 122373 208795 122439 208798
rect 68829 208178 68895 208181
rect 120717 208178 120783 208181
rect 68829 208176 70380 208178
rect 68829 208120 68834 208176
rect 68890 208120 70380 208176
rect 68829 208118 70380 208120
rect 119692 208176 120783 208178
rect 119692 208120 120722 208176
rect 120778 208120 120783 208176
rect 119692 208118 120783 208120
rect 68829 208115 68895 208118
rect 120717 208115 120783 208118
rect 167085 208178 167151 208181
rect 167085 208176 170292 208178
rect 167085 208120 167090 208176
rect 167146 208120 170292 208176
rect 167085 208118 170292 208120
rect 167085 208115 167151 208118
rect 69238 207436 69244 207500
rect 69308 207498 69314 207500
rect 230013 207498 230079 207501
rect 69308 207438 70380 207498
rect 229724 207496 230079 207498
rect 229724 207440 230018 207496
rect 230074 207440 230079 207496
rect 229724 207438 230079 207440
rect 69308 207436 69314 207438
rect 230013 207435 230079 207438
rect 121545 206818 121611 206821
rect 119692 206816 121611 206818
rect 3509 206274 3575 206277
rect 67725 206274 67791 206277
rect 70350 206274 70410 206788
rect 119692 206760 121550 206816
rect 121606 206760 121611 206816
rect 119692 206758 121611 206760
rect 121545 206755 121611 206758
rect 167085 206818 167151 206821
rect 168281 206818 168347 206821
rect 167085 206816 170292 206818
rect 167085 206760 167090 206816
rect 167146 206760 168286 206816
rect 168342 206760 170292 206816
rect 167085 206758 170292 206760
rect 167085 206755 167151 206758
rect 168281 206755 168347 206758
rect 3509 206272 70410 206274
rect 3509 206216 3514 206272
rect 3570 206216 67730 206272
rect 67786 206216 70410 206272
rect 3509 206214 70410 206216
rect 3509 206211 3575 206214
rect 67725 206211 67791 206214
rect 121545 206138 121611 206141
rect 119692 206136 121611 206138
rect 119692 206080 121550 206136
rect 121606 206080 121611 206136
rect 119692 206078 121611 206080
rect 121545 206075 121611 206078
rect 167085 206138 167151 206141
rect 167361 206138 167427 206141
rect 230657 206138 230723 206141
rect 232681 206138 232747 206141
rect 167085 206136 170292 206138
rect 167085 206080 167090 206136
rect 167146 206080 167366 206136
rect 167422 206080 170292 206136
rect 167085 206078 170292 206080
rect 229724 206136 232747 206138
rect 229724 206080 230662 206136
rect 230718 206080 232686 206136
rect 232742 206080 232747 206136
rect 229724 206078 232747 206080
rect 167085 206075 167151 206078
rect 167361 206075 167427 206078
rect 230657 206075 230723 206078
rect 232681 206075 232747 206078
rect 579981 205730 580047 205733
rect 583520 205730 584960 205820
rect 579981 205728 584960 205730
rect 579981 205672 579986 205728
rect 580042 205672 584960 205728
rect 579981 205670 584960 205672
rect 579981 205667 580047 205670
rect 67817 205594 67883 205597
rect 68502 205594 68508 205596
rect 67817 205592 68508 205594
rect 67817 205536 67822 205592
rect 67878 205536 68508 205592
rect 67817 205534 68508 205536
rect 67817 205531 67883 205534
rect 68502 205532 68508 205534
rect 68572 205594 68578 205596
rect 68572 205534 70380 205594
rect 583520 205580 584960 205670
rect 68572 205532 68578 205534
rect 121729 205458 121795 205461
rect 122557 205458 122623 205461
rect 119692 205456 122623 205458
rect 119692 205400 121734 205456
rect 121790 205400 122562 205456
rect 122618 205400 122623 205456
rect 119692 205398 122623 205400
rect 121729 205395 121795 205398
rect 122557 205395 122623 205398
rect 170121 205050 170187 205053
rect 170121 205048 170322 205050
rect 170121 204992 170126 205048
rect 170182 204992 170322 205048
rect 170121 204990 170322 204992
rect 170121 204987 170187 204990
rect 68921 204914 68987 204917
rect 69790 204914 69796 204916
rect 68921 204912 69796 204914
rect 68921 204856 68926 204912
rect 68982 204856 69796 204912
rect 68921 204854 69796 204856
rect 68921 204851 68987 204854
rect 69790 204852 69796 204854
rect 69860 204852 69866 204916
rect 68093 204778 68159 204781
rect 68093 204776 70380 204778
rect 68093 204720 68098 204776
rect 68154 204720 70380 204776
rect 68093 204718 70380 204720
rect 68093 204715 68159 204718
rect 167310 204716 167316 204780
rect 167380 204778 167386 204780
rect 170262 204778 170322 204990
rect 231894 204778 231900 204780
rect 167380 204748 170322 204778
rect 167380 204718 170292 204748
rect 229724 204718 231900 204778
rect 167380 204716 167386 204718
rect 231894 204716 231900 204718
rect 231964 204778 231970 204780
rect 233141 204778 233207 204781
rect 231964 204776 233207 204778
rect 231964 204720 233146 204776
rect 233202 204720 233207 204776
rect 231964 204718 233207 204720
rect 231964 204716 231970 204718
rect 233141 204715 233207 204718
rect 122557 204098 122623 204101
rect 229921 204098 229987 204101
rect 232681 204098 232747 204101
rect 119692 204096 122623 204098
rect 119692 204040 122562 204096
rect 122618 204040 122623 204096
rect 119692 204038 122623 204040
rect 229724 204096 232747 204098
rect 229724 204040 229926 204096
rect 229982 204040 232686 204096
rect 232742 204040 232747 204096
rect 229724 204038 232747 204040
rect 122557 204035 122623 204038
rect 229921 204035 229987 204038
rect 232681 204035 232747 204038
rect 68318 203356 68324 203420
rect 68388 203418 68394 203420
rect 120073 203418 120139 203421
rect 68388 203358 70380 203418
rect 119692 203416 120139 203418
rect 119692 203360 120078 203416
rect 120134 203360 120139 203416
rect 119692 203358 120139 203360
rect 68388 203356 68394 203358
rect 120073 203355 120139 203358
rect 167269 203418 167335 203421
rect 167269 203416 170292 203418
rect 167269 203360 167274 203416
rect 167330 203360 170292 203416
rect 167269 203358 170292 203360
rect 167269 203355 167335 203358
rect 229369 203010 229435 203013
rect 229326 203008 229435 203010
rect 229326 202952 229374 203008
rect 229430 202952 229435 203008
rect 229326 202947 229435 202952
rect 229326 202874 229386 202947
rect 229326 202814 229754 202874
rect 67633 202738 67699 202741
rect 167453 202738 167519 202741
rect 229694 202738 229754 202814
rect 232681 202738 232747 202741
rect 67633 202736 70380 202738
rect 67633 202680 67638 202736
rect 67694 202680 70380 202736
rect 67633 202678 70380 202680
rect 167453 202736 170292 202738
rect 167453 202680 167458 202736
rect 167514 202680 170292 202736
rect 229694 202736 232747 202738
rect 229694 202708 232686 202736
rect 167453 202678 170292 202680
rect 229724 202680 232686 202708
rect 232742 202680 232747 202736
rect 229724 202678 232747 202680
rect 67633 202675 67699 202678
rect 167453 202675 167519 202678
rect 232681 202675 232747 202678
rect 121821 202058 121887 202061
rect 119692 202056 121887 202058
rect -960 201922 480 202012
rect 119692 202000 121826 202056
rect 121882 202000 121887 202056
rect 119692 201998 121887 202000
rect 121821 201995 121887 201998
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 68645 201378 68711 201381
rect 120349 201378 120415 201381
rect 122557 201378 122623 201381
rect 68645 201376 70380 201378
rect 68645 201320 68650 201376
rect 68706 201320 70380 201376
rect 68645 201318 70380 201320
rect 119692 201376 122623 201378
rect 119692 201320 120354 201376
rect 120410 201320 122562 201376
rect 122618 201320 122623 201376
rect 119692 201318 122623 201320
rect 68645 201315 68711 201318
rect 120349 201315 120415 201318
rect 122557 201315 122623 201318
rect 167085 201378 167151 201381
rect 233325 201378 233391 201381
rect 167085 201376 170292 201378
rect 167085 201320 167090 201376
rect 167146 201320 170292 201376
rect 167085 201318 170292 201320
rect 229724 201376 233391 201378
rect 229724 201320 233330 201376
rect 233386 201320 233391 201376
rect 229724 201318 233391 201320
rect 167085 201315 167151 201318
rect 233325 201315 233391 201318
rect 68369 201242 68435 201245
rect 69606 201242 69612 201244
rect 68369 201240 69612 201242
rect 68369 201184 68374 201240
rect 68430 201184 69612 201240
rect 68369 201182 69612 201184
rect 68369 201179 68435 201182
rect 69606 201180 69612 201182
rect 69676 201180 69682 201244
rect 69289 200698 69355 200701
rect 232589 200698 232655 200701
rect 69289 200696 70380 200698
rect 69289 200640 69294 200696
rect 69350 200640 70380 200696
rect 69289 200638 70380 200640
rect 229724 200696 232655 200698
rect 229724 200640 232594 200696
rect 232650 200640 232655 200696
rect 229724 200638 232655 200640
rect 69289 200635 69355 200638
rect 232589 200635 232655 200638
rect 65425 200290 65491 200293
rect 70158 200290 70164 200292
rect 65425 200288 70164 200290
rect 65425 200232 65430 200288
rect 65486 200232 70164 200288
rect 65425 200230 70164 200232
rect 65425 200227 65491 200230
rect 70158 200228 70164 200230
rect 70228 200228 70234 200292
rect 70669 200290 70735 200293
rect 70534 200288 70735 200290
rect 70534 200232 70674 200288
rect 70730 200232 70735 200288
rect 70534 200230 70735 200232
rect 67398 200092 67404 200156
rect 67468 200154 67474 200156
rect 69238 200154 69244 200156
rect 67468 200094 69244 200154
rect 67468 200092 67474 200094
rect 69238 200092 69244 200094
rect 69308 200092 69314 200156
rect 70534 199885 70594 200230
rect 70669 200227 70735 200230
rect 167361 200018 167427 200021
rect 167361 200016 170292 200018
rect 70485 199880 70594 199885
rect 70485 199824 70490 199880
rect 70546 199824 70594 199880
rect 70485 199822 70594 199824
rect 70485 199819 70551 199822
rect 119662 199477 119722 199988
rect 167361 199960 167366 200016
rect 167422 199960 170292 200016
rect 167361 199958 170292 199960
rect 167361 199955 167427 199958
rect 119662 199472 119771 199477
rect 119662 199416 119710 199472
rect 119766 199416 119771 199472
rect 119662 199414 119771 199416
rect 119705 199411 119771 199414
rect 82077 199338 82143 199341
rect 84929 199338 84995 199341
rect 232681 199338 232747 199341
rect 82077 199336 84995 199338
rect 82077 199280 82082 199336
rect 82138 199280 84934 199336
rect 84990 199280 84995 199336
rect 82077 199278 84995 199280
rect 229724 199336 232747 199338
rect 229724 199280 232686 199336
rect 232742 199280 232747 199336
rect 229724 199278 232747 199280
rect 82077 199275 82143 199278
rect 84929 199275 84995 199278
rect 232681 199275 232747 199278
rect 68686 198732 68692 198796
rect 68756 198794 68762 198796
rect 72601 198794 72667 198797
rect 68756 198792 72667 198794
rect 68756 198736 72606 198792
rect 72662 198736 72667 198792
rect 68756 198734 72667 198736
rect 68756 198732 68762 198734
rect 72601 198731 72667 198734
rect 54477 198658 54543 198661
rect 107469 198658 107535 198661
rect 54477 198656 107535 198658
rect 54477 198600 54482 198656
rect 54538 198600 107474 198656
rect 107530 198600 107535 198656
rect 54477 198598 107535 198600
rect 54477 198595 54543 198598
rect 107469 198595 107535 198598
rect 103421 198522 103487 198525
rect 122833 198522 122899 198525
rect 103421 198520 122899 198522
rect 103421 198464 103426 198520
rect 103482 198464 122838 198520
rect 122894 198464 122899 198520
rect 103421 198462 122899 198464
rect 103421 198459 103487 198462
rect 122833 198459 122899 198462
rect 169886 198386 169892 198388
rect 161430 198326 169892 198386
rect 93853 198114 93919 198117
rect 161430 198114 161490 198326
rect 169886 198324 169892 198326
rect 169956 198324 169962 198388
rect 168925 198250 168991 198253
rect 170262 198250 170322 198628
rect 93853 198112 161490 198114
rect 93853 198056 93858 198112
rect 93914 198056 161490 198112
rect 93853 198054 161490 198056
rect 167134 198248 170322 198250
rect 167134 198192 168930 198248
rect 168986 198192 170322 198248
rect 167134 198190 170322 198192
rect 93853 198051 93919 198054
rect 66897 197978 66963 197981
rect 167134 197978 167194 198190
rect 168925 198187 168991 198190
rect 66897 197976 167194 197978
rect 66897 197920 66902 197976
rect 66958 197920 167194 197976
rect 66897 197918 167194 197920
rect 167361 197978 167427 197981
rect 232589 197978 232655 197981
rect 167361 197976 170292 197978
rect 167361 197920 167366 197976
rect 167422 197920 170292 197976
rect 167361 197918 170292 197920
rect 229724 197976 232655 197978
rect 229724 197920 232594 197976
rect 232650 197920 232655 197976
rect 229724 197918 232655 197920
rect 66897 197915 66963 197918
rect 167361 197915 167427 197918
rect 232589 197915 232655 197918
rect 108849 196754 108915 196757
rect 119286 196754 119292 196756
rect 108849 196752 119292 196754
rect 108849 196696 108854 196752
rect 108910 196696 119292 196752
rect 108849 196694 119292 196696
rect 108849 196691 108915 196694
rect 119286 196692 119292 196694
rect 119356 196692 119362 196756
rect 108573 196618 108639 196621
rect 120206 196618 120212 196620
rect 108573 196616 120212 196618
rect 108573 196560 108578 196616
rect 108634 196560 120212 196616
rect 108573 196558 120212 196560
rect 108573 196555 108639 196558
rect 120206 196556 120212 196558
rect 120276 196556 120282 196620
rect 167361 196618 167427 196621
rect 167361 196616 170292 196618
rect 167361 196560 167366 196616
rect 167422 196560 170292 196616
rect 167361 196558 170292 196560
rect 167361 196555 167427 196558
rect 229326 196213 229386 196588
rect 229326 196208 229435 196213
rect 229326 196152 229374 196208
rect 229430 196152 229435 196208
rect 229326 196150 229435 196152
rect 229369 196147 229435 196150
rect 229510 195397 229570 195908
rect 229461 195392 229570 195397
rect 229461 195336 229466 195392
rect 229522 195336 229570 195392
rect 229461 195334 229570 195336
rect 229461 195331 229527 195334
rect 167678 195196 167684 195260
rect 167748 195258 167754 195260
rect 168189 195258 168255 195261
rect 167748 195256 170292 195258
rect 167748 195200 168194 195256
rect 168250 195200 170292 195256
rect 167748 195198 170292 195200
rect 167748 195196 167754 195198
rect 168189 195195 168255 195198
rect 69790 194516 69796 194580
rect 69860 194578 69866 194580
rect 169937 194578 170003 194581
rect 232405 194578 232471 194581
rect 69860 194576 170292 194578
rect 69860 194520 169942 194576
rect 169998 194520 170292 194576
rect 69860 194518 170292 194520
rect 229724 194576 232471 194578
rect 229724 194520 232410 194576
rect 232466 194520 232471 194576
rect 229724 194518 232471 194520
rect 69860 194516 69866 194518
rect 169937 194515 170003 194518
rect 232405 194515 232471 194518
rect 167862 193156 167868 193220
rect 167932 193218 167938 193220
rect 168281 193218 168347 193221
rect 167932 193216 170292 193218
rect 167932 193160 168286 193216
rect 168342 193160 170292 193216
rect 167932 193158 170292 193160
rect 167932 193156 167938 193158
rect 168281 193155 168347 193158
rect 229510 192813 229570 193188
rect 229510 192808 229619 192813
rect 229510 192752 229558 192808
rect 229614 192752 229619 192808
rect 229510 192750 229619 192752
rect 229553 192747 229619 192750
rect 112989 192538 113055 192541
rect 122230 192538 122236 192540
rect 112989 192536 122236 192538
rect 112989 192480 112994 192536
rect 113050 192480 122236 192536
rect 112989 192478 122236 192480
rect 112989 192475 113055 192478
rect 122230 192476 122236 192478
rect 122300 192476 122306 192540
rect 232313 192538 232379 192541
rect 229724 192536 232379 192538
rect 229724 192480 232318 192536
rect 232374 192480 232379 192536
rect 229724 192478 232379 192480
rect 232313 192475 232379 192478
rect 579705 192538 579771 192541
rect 583520 192538 584960 192628
rect 579705 192536 584960 192538
rect 579705 192480 579710 192536
rect 579766 192480 584960 192536
rect 579705 192478 584960 192480
rect 579705 192475 579771 192478
rect 583520 192388 584960 192478
rect 167361 191858 167427 191861
rect 167361 191856 170292 191858
rect 167361 191800 167366 191856
rect 167422 191800 170292 191856
rect 167361 191798 170292 191800
rect 167361 191795 167427 191798
rect 233141 191178 233207 191181
rect 229724 191176 233207 191178
rect 229724 191120 233146 191176
rect 233202 191120 233207 191176
rect 229724 191118 233207 191120
rect 233141 191115 233207 191118
rect 168097 190498 168163 190501
rect 169569 190498 169635 190501
rect 168097 190496 170292 190498
rect 168097 190440 168102 190496
rect 168158 190440 169574 190496
rect 169630 190440 170292 190496
rect 168097 190438 170292 190440
rect 168097 190435 168163 190438
rect 169569 190435 169635 190438
rect 167361 189818 167427 189821
rect 232221 189818 232287 189821
rect 167361 189816 170292 189818
rect 167361 189760 167366 189816
rect 167422 189760 170292 189816
rect 167361 189758 170292 189760
rect 229724 189816 232287 189818
rect 229724 189760 232226 189816
rect 232282 189760 232287 189816
rect 229724 189758 232287 189760
rect 167361 189755 167427 189758
rect 232221 189755 232287 189758
rect -960 188866 480 188956
rect 69606 188940 69612 189004
rect 69676 189002 69682 189004
rect 169845 189002 169911 189005
rect 69676 189000 170322 189002
rect 69676 188944 169850 189000
rect 169906 188944 170322 189000
rect 69676 188942 170322 188944
rect 69676 188940 69682 188942
rect 169845 188939 169911 188942
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 170262 188428 170322 188942
rect 232773 188458 232839 188461
rect 229724 188456 232839 188458
rect 229724 188400 232778 188456
rect 232834 188400 232839 188456
rect 229724 188398 232839 188400
rect 232773 188395 232839 188398
rect 233141 187778 233207 187781
rect 229724 187776 233207 187778
rect 229724 187720 233146 187776
rect 233202 187720 233207 187776
rect 229724 187718 233207 187720
rect 233141 187715 233207 187718
rect 68185 186690 68251 186693
rect 170262 186690 170322 187068
rect 68185 186688 170322 186690
rect 68185 186632 68190 186688
rect 68246 186632 170322 186688
rect 68185 186630 170322 186632
rect 68185 186627 68251 186630
rect 167361 186418 167427 186421
rect 233141 186418 233207 186421
rect 167361 186416 170292 186418
rect 167361 186360 167366 186416
rect 167422 186360 170292 186416
rect 167361 186358 170292 186360
rect 229724 186416 233207 186418
rect 229724 186360 233146 186416
rect 233202 186360 233207 186416
rect 229724 186358 233207 186360
rect 167361 186355 167427 186358
rect 233141 186355 233207 186358
rect 167361 185058 167427 185061
rect 168281 185058 168347 185061
rect 231853 185058 231919 185061
rect 167361 185056 170292 185058
rect 167361 185000 167366 185056
rect 167422 185000 168286 185056
rect 168342 185000 170292 185056
rect 167361 184998 170292 185000
rect 229724 185056 231919 185058
rect 229724 185000 231858 185056
rect 231914 185000 231919 185056
rect 229724 184998 231919 185000
rect 167361 184995 167427 184998
rect 168281 184995 168347 184998
rect 231853 184995 231919 184998
rect 232129 184378 232195 184381
rect 229724 184376 232195 184378
rect 229724 184320 232134 184376
rect 232190 184320 232195 184376
rect 229724 184318 232195 184320
rect 232129 184315 232195 184318
rect 167361 183698 167427 183701
rect 167361 183696 170292 183698
rect 167361 183640 167366 183696
rect 167422 183640 170292 183696
rect 167361 183638 170292 183640
rect 167361 183635 167427 183638
rect 232405 183018 232471 183021
rect 229724 183016 232471 183018
rect 229724 182960 232410 183016
rect 232466 182960 232471 183016
rect 229724 182958 232471 182960
rect 232405 182955 232471 182958
rect 167361 182338 167427 182341
rect 167361 182336 170292 182338
rect 167361 182280 167366 182336
rect 167422 182280 170292 182336
rect 167361 182278 170292 182280
rect 167361 182275 167427 182278
rect 67725 180978 67791 180981
rect 71262 180978 71268 180980
rect 67725 180976 71268 180978
rect 67725 180920 67730 180976
rect 67786 180920 71268 180976
rect 67725 180918 71268 180920
rect 67725 180915 67791 180918
rect 71262 180916 71268 180918
rect 71332 180916 71338 180980
rect 71078 180780 71084 180844
rect 71148 180842 71154 180844
rect 170262 180842 170322 181628
rect 229694 181117 229754 181628
rect 229694 181112 229803 181117
rect 229694 181056 229742 181112
rect 229798 181056 229803 181112
rect 229694 181054 229803 181056
rect 229737 181051 229803 181054
rect 71148 180782 170322 180842
rect 71148 180780 71154 180782
rect 167453 180298 167519 180301
rect 168189 180298 168255 180301
rect 232221 180298 232287 180301
rect 167453 180296 170292 180298
rect 167453 180240 167458 180296
rect 167514 180240 168194 180296
rect 168250 180240 170292 180296
rect 167453 180238 170292 180240
rect 229724 180296 232287 180298
rect 229724 180240 232226 180296
rect 232282 180240 232287 180296
rect 229724 180238 232287 180240
rect 167453 180235 167519 180238
rect 168189 180235 168255 180238
rect 232221 180235 232287 180238
rect 231853 179618 231919 179621
rect 229724 179616 231919 179618
rect 229724 179560 231858 179616
rect 231914 179560 231919 179616
rect 229724 179558 231919 179560
rect 231853 179555 231919 179558
rect 69238 179284 69244 179348
rect 69308 179346 69314 179348
rect 169661 179346 169727 179349
rect 69308 179344 170322 179346
rect 69308 179288 169666 179344
rect 169722 179288 170322 179344
rect 69308 179286 170322 179288
rect 69308 179284 69314 179286
rect 169661 179283 169727 179286
rect 170262 178908 170322 179286
rect 580257 179210 580323 179213
rect 583520 179210 584960 179300
rect 580257 179208 584960 179210
rect 580257 179152 580262 179208
rect 580318 179152 584960 179208
rect 580257 179150 584960 179152
rect 580257 179147 580323 179150
rect 583520 179060 584960 179150
rect 232037 178258 232103 178261
rect 229724 178256 232103 178258
rect 71262 178060 71268 178124
rect 71332 178122 71338 178124
rect 170262 178122 170322 178228
rect 229724 178200 232042 178256
rect 232098 178200 232103 178256
rect 229724 178198 232103 178200
rect 232037 178195 232103 178198
rect 71332 178062 170322 178122
rect 71332 178060 71338 178062
rect 68502 177244 68508 177308
rect 68572 177306 68578 177308
rect 68921 177306 68987 177309
rect 68572 177304 68987 177306
rect 68572 177248 68926 177304
rect 68982 177248 68987 177304
rect 68572 177246 68987 177248
rect 68572 177244 68578 177246
rect 68921 177243 68987 177246
rect 167453 176898 167519 176901
rect 232497 176898 232563 176901
rect 167453 176896 170292 176898
rect 167453 176840 167458 176896
rect 167514 176840 170292 176896
rect 167453 176838 170292 176840
rect 229724 176896 232563 176898
rect 229724 176840 232502 176896
rect 232558 176840 232563 176896
rect 229724 176838 232563 176840
rect 167453 176835 167519 176838
rect 232497 176835 232563 176838
rect 231945 176218 232011 176221
rect 229724 176216 232011 176218
rect 229724 176160 231950 176216
rect 232006 176160 232011 176216
rect 229724 176158 232011 176160
rect 231945 176155 232011 176158
rect -960 175796 480 176036
rect 69238 175884 69244 175948
rect 69308 175946 69314 175948
rect 69381 175946 69447 175949
rect 69308 175944 69447 175946
rect 69308 175888 69386 175944
rect 69442 175888 69447 175944
rect 69308 175886 69447 175888
rect 69308 175884 69314 175886
rect 69381 175883 69447 175886
rect 112897 175946 112963 175949
rect 122414 175946 122420 175948
rect 112897 175944 122420 175946
rect 112897 175888 112902 175944
rect 112958 175888 122420 175944
rect 112897 175886 122420 175888
rect 112897 175883 112963 175886
rect 122414 175884 122420 175886
rect 122484 175884 122490 175948
rect 168097 175538 168163 175541
rect 169518 175538 169524 175540
rect 168097 175536 169524 175538
rect 168097 175480 168102 175536
rect 168158 175480 169524 175536
rect 168097 175478 169524 175480
rect 168097 175475 168163 175478
rect 169518 175476 169524 175478
rect 169588 175538 169594 175540
rect 169588 175478 170292 175538
rect 169588 175476 169594 175478
rect 231025 174858 231091 174861
rect 233049 174858 233115 174861
rect 229724 174856 233115 174858
rect 229724 174800 231030 174856
rect 231086 174800 233054 174856
rect 233110 174800 233115 174856
rect 229724 174798 233115 174800
rect 231025 174795 231091 174798
rect 233049 174795 233115 174798
rect 68318 173980 68324 174044
rect 68388 174042 68394 174044
rect 170262 174042 170322 174148
rect 68388 173982 170322 174042
rect 68388 173980 68394 173982
rect 168741 173498 168807 173501
rect 169109 173498 169175 173501
rect 232037 173498 232103 173501
rect 168741 173496 170292 173498
rect 168741 173440 168746 173496
rect 168802 173440 169114 173496
rect 169170 173440 170292 173496
rect 168741 173438 170292 173440
rect 229724 173496 232103 173498
rect 229724 173440 232042 173496
rect 232098 173440 232103 173496
rect 229724 173438 232103 173440
rect 168741 173435 168807 173438
rect 169109 173435 169175 173438
rect 232037 173435 232103 173438
rect 168097 172138 168163 172141
rect 168097 172136 170292 172138
rect 168097 172080 168102 172136
rect 168158 172080 170292 172136
rect 168097 172078 170292 172080
rect 168097 172075 168163 172078
rect 229694 171866 229754 172108
rect 231761 171866 231827 171869
rect 229694 171864 231827 171866
rect 229694 171808 231766 171864
rect 231822 171808 231827 171864
rect 229694 171806 231827 171808
rect 231761 171803 231827 171806
rect 229694 171186 229754 171428
rect 231669 171186 231735 171189
rect 229694 171184 231735 171186
rect 229694 171128 231674 171184
rect 231730 171128 231735 171184
rect 229694 171126 231735 171128
rect 231669 171123 231735 171126
rect 168097 170778 168163 170781
rect 168097 170776 170292 170778
rect 168097 170720 168102 170776
rect 168158 170720 170292 170776
rect 168097 170718 170292 170720
rect 168097 170715 168163 170718
rect 233877 170098 233943 170101
rect 229540 170096 233943 170098
rect 229540 170068 233882 170096
rect 229510 170040 233882 170068
rect 233938 170040 233943 170096
rect 229510 170038 233943 170040
rect 170305 169690 170371 169693
rect 221549 169690 221615 169693
rect 170305 169688 221615 169690
rect 170305 169632 170310 169688
rect 170366 169632 221554 169688
rect 221610 169632 221615 169688
rect 170305 169630 221615 169632
rect 170305 169627 170371 169630
rect 221549 169627 221615 169630
rect 165429 169554 165495 169557
rect 169886 169554 169892 169556
rect 165429 169552 169892 169554
rect 165429 169496 165434 169552
rect 165490 169496 169892 169552
rect 165429 169494 169892 169496
rect 165429 169491 165495 169494
rect 169886 169492 169892 169494
rect 169956 169554 169962 169556
rect 198365 169554 198431 169557
rect 169956 169552 198431 169554
rect 169956 169496 198370 169552
rect 198426 169496 198431 169552
rect 169956 169494 198431 169496
rect 169956 169492 169962 169494
rect 198365 169491 198431 169494
rect 229277 169554 229343 169557
rect 229510 169554 229570 170038
rect 233877 170035 233943 170038
rect 229277 169552 229570 169554
rect 229277 169496 229282 169552
rect 229338 169496 229570 169552
rect 229277 169494 229570 169496
rect 229277 169491 229343 169494
rect 74533 169010 74599 169013
rect 107009 169010 107075 169013
rect 175181 169010 175247 169013
rect 74533 169008 175247 169010
rect 74533 168952 74538 169008
rect 74594 168952 107014 169008
rect 107070 168952 175186 169008
rect 175242 168952 175247 169008
rect 74533 168950 175247 168952
rect 74533 168947 74599 168950
rect 107009 168947 107075 168950
rect 175181 168947 175247 168950
rect 170949 168330 171015 168333
rect 184933 168330 184999 168333
rect 170949 168328 184999 168330
rect 170949 168272 170954 168328
rect 171010 168272 184938 168328
rect 184994 168272 184999 168328
rect 170949 168270 184999 168272
rect 170949 168267 171015 168270
rect 184933 168267 184999 168270
rect 199326 168268 199332 168332
rect 199396 168330 199402 168332
rect 199653 168330 199719 168333
rect 199396 168328 199719 168330
rect 199396 168272 199658 168328
rect 199714 168272 199719 168328
rect 199396 168270 199719 168272
rect 199396 168268 199402 168270
rect 199653 168267 199719 168270
rect 168925 168194 168991 168197
rect 218329 168194 218395 168197
rect 168925 168192 218395 168194
rect 168925 168136 168930 168192
rect 168986 168136 218334 168192
rect 218390 168136 218395 168192
rect 168925 168134 218395 168136
rect 168925 168131 168991 168134
rect 218329 168131 218395 168134
rect 164877 168058 164943 168061
rect 193213 168058 193279 168061
rect 164877 168056 193279 168058
rect 164877 168000 164882 168056
rect 164938 168000 193218 168056
rect 193274 168000 193279 168056
rect 164877 167998 193279 168000
rect 164877 167995 164943 167998
rect 193213 167995 193279 167998
rect 168741 167922 168807 167925
rect 182909 167922 182975 167925
rect 168741 167920 182975 167922
rect 168741 167864 168746 167920
rect 168802 167864 182914 167920
rect 182970 167864 182975 167920
rect 168741 167862 182975 167864
rect 168741 167859 168807 167862
rect 182909 167859 182975 167862
rect 166533 167786 166599 167789
rect 226057 167786 226123 167789
rect 166533 167784 226123 167786
rect 166533 167728 166538 167784
rect 166594 167728 226062 167784
rect 226118 167728 226123 167784
rect 166533 167726 226123 167728
rect 166533 167723 166599 167726
rect 226057 167723 226123 167726
rect 120625 166972 120691 166973
rect 120574 166970 120580 166972
rect 120498 166910 120580 166970
rect 120644 166970 120691 166972
rect 233325 166970 233391 166973
rect 120644 166968 233391 166970
rect 120686 166912 233330 166968
rect 233386 166912 233391 166968
rect 120574 166908 120580 166910
rect 120644 166910 233391 166912
rect 120644 166908 120691 166910
rect 120625 166907 120691 166908
rect 233325 166907 233391 166910
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect 119102 165548 119108 165612
rect 119172 165610 119178 165612
rect 119337 165610 119403 165613
rect 119172 165608 119403 165610
rect 119172 165552 119342 165608
rect 119398 165552 119403 165608
rect 119172 165550 119403 165552
rect 119172 165548 119178 165550
rect 119337 165547 119403 165550
rect 156781 165610 156847 165613
rect 233601 165610 233667 165613
rect 156781 165608 233667 165610
rect 156781 165552 156786 165608
rect 156842 165552 233606 165608
rect 233662 165552 233667 165608
rect 156781 165550 233667 165552
rect 156781 165547 156847 165550
rect 233601 165547 233667 165550
rect -960 162890 480 162980
rect 3417 162890 3483 162893
rect -960 162888 3483 162890
rect -960 162832 3422 162888
rect 3478 162832 3483 162888
rect -960 162830 3483 162832
rect -960 162740 480 162830
rect 3417 162827 3483 162830
rect 580257 152690 580323 152693
rect 583520 152690 584960 152780
rect 580257 152688 584960 152690
rect 580257 152632 580262 152688
rect 580318 152632 584960 152688
rect 580257 152630 584960 152632
rect 580257 152627 580323 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 2957 149834 3023 149837
rect -960 149832 3023 149834
rect -960 149776 2962 149832
rect 3018 149776 3023 149832
rect -960 149774 3023 149776
rect -960 149684 480 149774
rect 2957 149771 3023 149774
rect 580257 139362 580323 139365
rect 583520 139362 584960 139452
rect 580257 139360 584960 139362
rect 580257 139304 580262 139360
rect 580318 139304 584960 139360
rect 580257 139302 584960 139304
rect 580257 139299 580323 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 119245 125490 119311 125493
rect 119654 125490 119660 125492
rect 119245 125488 119660 125490
rect 119245 125432 119250 125488
rect 119306 125432 119660 125488
rect 119245 125430 119660 125432
rect 119245 125427 119311 125430
rect 119654 125428 119660 125430
rect 119724 125428 119730 125492
rect 118918 125292 118924 125356
rect 118988 125354 118994 125356
rect 119705 125354 119771 125357
rect 118988 125352 119771 125354
rect 118988 125296 119710 125352
rect 119766 125296 119771 125352
rect 118988 125294 119771 125296
rect 118988 125292 118994 125294
rect 119705 125291 119771 125294
rect 117037 124538 117103 124541
rect 117037 124536 122850 124538
rect 117037 124480 117042 124536
rect 117098 124480 122850 124536
rect 117037 124478 122850 124480
rect 117037 124475 117103 124478
rect 122790 124266 122850 124478
rect 199510 124266 199516 124268
rect 122790 124206 199516 124266
rect 199510 124204 199516 124206
rect 199580 124204 199586 124268
rect -960 123572 480 123812
rect 111517 123450 111583 123453
rect 121862 123450 121868 123452
rect 111517 123448 121868 123450
rect 111517 123392 111522 123448
rect 111578 123392 121868 123448
rect 111517 123390 121868 123392
rect 111517 123387 111583 123390
rect 121862 123388 121868 123390
rect 121932 123388 121938 123452
rect 122046 122844 122052 122908
rect 122116 122906 122122 122908
rect 122189 122906 122255 122909
rect 204437 122906 204503 122909
rect 122116 122904 204503 122906
rect 122116 122848 122194 122904
rect 122250 122848 204442 122904
rect 204498 122848 204503 122904
rect 122116 122846 204503 122848
rect 122116 122844 122122 122846
rect 122189 122843 122255 122846
rect 204437 122843 204503 122846
rect 165981 122226 166047 122229
rect 191281 122226 191347 122229
rect 165981 122224 191347 122226
rect 165981 122168 165986 122224
rect 166042 122168 191286 122224
rect 191342 122168 191347 122224
rect 165981 122166 191347 122168
rect 165981 122163 166047 122166
rect 191281 122163 191347 122166
rect 164141 122090 164207 122093
rect 186773 122090 186839 122093
rect 164141 122088 186839 122090
rect 164141 122032 164146 122088
rect 164202 122032 186778 122088
rect 186834 122032 186839 122088
rect 164141 122030 186839 122032
rect 164141 122027 164207 122030
rect 186773 122027 186839 122030
rect 166533 121954 166599 121957
rect 178401 121954 178467 121957
rect 166533 121952 178467 121954
rect 166533 121896 166538 121952
rect 166594 121896 178406 121952
rect 178462 121896 178467 121952
rect 166533 121894 178467 121896
rect 166533 121891 166599 121894
rect 178401 121891 178467 121894
rect 168649 121818 168715 121821
rect 192569 121818 192635 121821
rect 168649 121816 192635 121818
rect 168649 121760 168654 121816
rect 168710 121760 192574 121816
rect 192630 121760 192635 121816
rect 168649 121758 192635 121760
rect 168649 121755 168715 121758
rect 192569 121755 192635 121758
rect 169937 121682 170003 121685
rect 180977 121682 181043 121685
rect 169937 121680 181043 121682
rect 169937 121624 169942 121680
rect 169998 121624 180982 121680
rect 181038 121624 181043 121680
rect 169937 121622 181043 121624
rect 169937 121619 170003 121622
rect 180977 121619 181043 121622
rect 131113 121410 131179 121413
rect 131849 121410 131915 121413
rect 193121 121410 193187 121413
rect 131113 121408 193187 121410
rect 131113 121352 131118 121408
rect 131174 121352 131854 121408
rect 131910 121352 193126 121408
rect 193182 121352 193187 121408
rect 131113 121350 193187 121352
rect 131113 121347 131179 121350
rect 131849 121347 131915 121350
rect 193121 121347 193187 121350
rect 170070 120668 170076 120732
rect 170140 120730 170146 120732
rect 193213 120730 193279 120733
rect 170140 120728 193279 120730
rect 170140 120672 193218 120728
rect 193274 120672 193279 120728
rect 170140 120670 193279 120672
rect 170140 120668 170146 120670
rect 193213 120667 193279 120670
rect 168465 120594 168531 120597
rect 180333 120594 180399 120597
rect 168465 120592 180399 120594
rect 168465 120536 168470 120592
rect 168526 120536 180338 120592
rect 180394 120536 180399 120592
rect 168465 120534 180399 120536
rect 168465 120531 168531 120534
rect 180333 120531 180399 120534
rect 169886 120396 169892 120460
rect 169956 120458 169962 120460
rect 182265 120458 182331 120461
rect 169956 120456 182331 120458
rect 169956 120400 182270 120456
rect 182326 120400 182331 120456
rect 169956 120398 182331 120400
rect 169956 120396 169962 120398
rect 182265 120395 182331 120398
rect 168373 120322 168439 120325
rect 188705 120322 188771 120325
rect 168373 120320 188771 120322
rect 168373 120264 168378 120320
rect 168434 120264 188710 120320
rect 188766 120264 188771 120320
rect 168373 120262 188771 120264
rect 168373 120259 168439 120262
rect 188705 120259 188771 120262
rect 169702 120124 169708 120188
rect 169772 120186 169778 120188
rect 175181 120186 175247 120189
rect 169772 120184 175247 120186
rect 169772 120128 175186 120184
rect 175242 120128 175247 120184
rect 169772 120126 175247 120128
rect 169772 120124 169778 120126
rect 175181 120123 175247 120126
rect 166901 119642 166967 119645
rect 166901 119640 170292 119642
rect 166901 119584 166906 119640
rect 166962 119584 170292 119640
rect 166901 119582 170292 119584
rect 166901 119579 166967 119582
rect 166022 119308 166028 119372
rect 166092 119370 166098 119372
rect 170673 119370 170739 119373
rect 200113 119372 200179 119373
rect 166092 119368 170739 119370
rect 166092 119312 170678 119368
rect 170734 119312 170739 119368
rect 166092 119310 170739 119312
rect 166092 119308 166098 119310
rect 170673 119307 170739 119310
rect 200062 119308 200068 119372
rect 200132 119370 200179 119372
rect 200132 119368 200224 119370
rect 200174 119312 200224 119368
rect 200132 119310 200224 119312
rect 200132 119308 200179 119310
rect 200113 119307 200179 119308
rect 199694 119036 199700 119100
rect 199764 119036 199770 119100
rect 166942 118764 166948 118828
rect 167012 118826 167018 118828
rect 167269 118826 167335 118829
rect 167012 118824 167335 118826
rect 167012 118768 167274 118824
rect 167330 118768 167335 118824
rect 167012 118766 167335 118768
rect 167012 118764 167018 118766
rect 167269 118763 167335 118766
rect 200062 118628 200068 118692
rect 200132 118690 200138 118692
rect 201953 118690 202019 118693
rect 200132 118688 202019 118690
rect 200132 118632 201958 118688
rect 202014 118632 202019 118688
rect 200132 118630 202019 118632
rect 200132 118628 200138 118630
rect 201953 118627 202019 118630
rect 199694 118356 199700 118420
rect 199764 118356 199770 118420
rect 167085 118282 167151 118285
rect 169201 118282 169267 118285
rect 167085 118280 170292 118282
rect 167085 118224 167090 118280
rect 167146 118224 169206 118280
rect 169262 118224 170292 118280
rect 167085 118222 170292 118224
rect 167085 118219 167151 118222
rect 169201 118219 169267 118222
rect 76465 118010 76531 118013
rect 166022 118010 166028 118012
rect 76465 118008 166028 118010
rect 76465 117952 76470 118008
rect 76526 117952 166028 118008
rect 76465 117950 166028 117952
rect 76465 117947 76531 117950
rect 166022 117948 166028 117950
rect 166092 117948 166098 118012
rect 200062 117948 200068 118012
rect 200132 118010 200138 118012
rect 201953 118010 202019 118013
rect 200132 118008 202019 118010
rect 200132 117952 201958 118008
rect 202014 117952 202019 118008
rect 200132 117950 202019 117952
rect 200132 117948 200138 117950
rect 201953 117947 202019 117950
rect 199694 117676 199700 117740
rect 199764 117676 199770 117740
rect 166993 117602 167059 117605
rect 166993 117600 170292 117602
rect 166993 117544 166998 117600
rect 167054 117544 170292 117600
rect 166993 117542 170292 117544
rect 166993 117539 167059 117542
rect 68829 117332 68895 117333
rect 68829 117330 68876 117332
rect 68784 117328 68876 117330
rect 68784 117272 68834 117328
rect 68784 117270 68876 117272
rect 68829 117268 68876 117270
rect 68940 117268 68946 117332
rect 200062 117268 200068 117332
rect 200132 117330 200138 117332
rect 202137 117330 202203 117333
rect 200132 117328 202203 117330
rect 200132 117272 202142 117328
rect 202198 117272 202203 117328
rect 200132 117270 202203 117272
rect 200132 117268 200138 117270
rect 68829 117267 68895 117268
rect 202137 117267 202203 117270
rect 199694 116996 199700 117060
rect 199764 116996 199770 117060
rect 170254 116860 170260 116924
rect 170324 116860 170330 116924
rect 170262 116650 170322 116860
rect 170078 116590 170322 116650
rect 76465 116514 76531 116517
rect 166942 116514 166948 116516
rect 76465 116512 166948 116514
rect 76465 116456 76470 116512
rect 76526 116456 166948 116512
rect 76465 116454 166948 116456
rect 76465 116451 76531 116454
rect 166942 116452 166948 116454
rect 167012 116452 167018 116516
rect 73245 116242 73311 116245
rect 170078 116242 170138 116590
rect 199510 116316 199516 116380
rect 199580 116316 199586 116380
rect 73245 116240 170138 116242
rect 73245 116184 73250 116240
rect 73306 116184 170138 116240
rect 73245 116182 170138 116184
rect 73245 116179 73311 116182
rect 68829 116106 68895 116109
rect 168925 116106 168991 116109
rect 68829 116104 168991 116106
rect 68829 116048 68834 116104
rect 68890 116048 168930 116104
rect 168986 116048 168991 116104
rect 68829 116046 168991 116048
rect 68829 116043 68895 116046
rect 168925 116043 168991 116046
rect 169109 116106 169175 116109
rect 169569 116106 169635 116109
rect 170262 116106 170322 116212
rect 169109 116104 170322 116106
rect 169109 116048 169114 116104
rect 169170 116048 169574 116104
rect 169630 116048 170322 116104
rect 169109 116046 170322 116048
rect 169109 116043 169175 116046
rect 169569 116043 169635 116046
rect 200062 115908 200068 115972
rect 200132 115908 200138 115972
rect 200070 115834 200130 115908
rect 202413 115834 202479 115837
rect 200070 115832 202479 115834
rect 200070 115776 202418 115832
rect 202474 115776 202479 115832
rect 200070 115774 202479 115776
rect 202413 115771 202479 115774
rect 199694 115636 199700 115700
rect 199764 115636 199770 115700
rect 166993 115562 167059 115565
rect 166993 115560 170292 115562
rect 166993 115504 166998 115560
rect 167054 115504 170292 115560
rect 166993 115502 170292 115504
rect 166993 115499 167059 115502
rect 200062 115228 200068 115292
rect 200132 115290 200138 115292
rect 201953 115290 202019 115293
rect 200132 115288 202019 115290
rect 200132 115232 201958 115288
rect 202014 115232 202019 115288
rect 200132 115230 202019 115232
rect 200132 115228 200138 115230
rect 201953 115227 202019 115230
rect 199694 114956 199700 115020
rect 199764 114956 199770 115020
rect 167177 114882 167243 114885
rect 170254 114882 170260 114884
rect 167177 114880 170260 114882
rect 167177 114824 167182 114880
rect 167238 114824 170260 114880
rect 167177 114822 170260 114824
rect 167177 114819 167243 114822
rect 170254 114820 170260 114822
rect 170324 114820 170330 114884
rect 200062 114548 200068 114612
rect 200132 114548 200138 114612
rect 200070 114474 200130 114548
rect 202321 114474 202387 114477
rect 200070 114472 202387 114474
rect 200070 114416 202326 114472
rect 202382 114416 202387 114472
rect 200070 114414 202387 114416
rect 202321 114411 202387 114414
rect 169293 114202 169359 114205
rect 169293 114200 170292 114202
rect 169293 114144 169298 114200
rect 169354 114144 170292 114200
rect 169293 114142 170292 114144
rect 169293 114139 169359 114142
rect 143441 114066 143507 114069
rect 170070 114066 170076 114068
rect 143441 114064 170076 114066
rect 143441 114008 143446 114064
rect 143502 114008 170076 114064
rect 143441 114006 170076 114008
rect 143441 114003 143507 114006
rect 170070 114004 170076 114006
rect 170140 114004 170146 114068
rect 153009 113930 153075 113933
rect 169886 113930 169892 113932
rect 153009 113928 169892 113930
rect 153009 113872 153014 113928
rect 153070 113872 169892 113928
rect 153009 113870 169892 113872
rect 153009 113867 153075 113870
rect 169886 113868 169892 113870
rect 169956 113868 169962 113932
rect 140773 113794 140839 113797
rect 141417 113794 141483 113797
rect 169702 113794 169708 113796
rect 140773 113792 169708 113794
rect 140773 113736 140778 113792
rect 140834 113736 141422 113792
rect 141478 113736 169708 113792
rect 140773 113734 169708 113736
rect 140773 113731 140839 113734
rect 141417 113731 141483 113734
rect 169702 113732 169708 113734
rect 169772 113732 169778 113796
rect 199694 113596 199700 113660
rect 199764 113596 199770 113660
rect 200062 113188 200068 113252
rect 200132 113250 200138 113252
rect 200132 113190 200498 113250
rect 200132 113188 200138 113190
rect 200113 113114 200179 113117
rect 200070 113112 200179 113114
rect 200070 113056 200118 113112
rect 200174 113056 200179 113112
rect 200070 113051 200179 113056
rect 200297 113114 200363 113117
rect 200438 113114 200498 113190
rect 200297 113112 200498 113114
rect 200297 113056 200302 113112
rect 200358 113056 200498 113112
rect 200297 113054 200498 113056
rect 200297 113051 200363 113054
rect 169385 112842 169451 112845
rect 169385 112840 170292 112842
rect 169385 112784 169390 112840
rect 169446 112784 170292 112840
rect 169385 112782 170292 112784
rect 169385 112779 169451 112782
rect 199694 112780 199700 112844
rect 199764 112780 199770 112844
rect 200070 112572 200130 113051
rect 580349 112842 580415 112845
rect 583520 112842 584960 112932
rect 580349 112840 584960 112842
rect 580349 112784 580354 112840
rect 580410 112784 584960 112840
rect 580349 112782 584960 112784
rect 580349 112779 580415 112782
rect 583520 112692 584960 112782
rect 70526 112508 70532 112572
rect 70596 112570 70602 112572
rect 70596 112510 80070 112570
rect 70596 112508 70602 112510
rect 67214 112372 67220 112436
rect 67284 112434 67290 112436
rect 67284 112374 75194 112434
rect 67284 112372 67290 112374
rect 66069 112162 66135 112165
rect 74993 112162 75059 112165
rect 66069 112160 75059 112162
rect 66069 112104 66074 112160
rect 66130 112104 74998 112160
rect 75054 112104 75059 112160
rect 66069 112102 75059 112104
rect 75134 112162 75194 112374
rect 80010 112298 80070 112510
rect 200062 112508 200068 112572
rect 200132 112508 200138 112572
rect 150433 112298 150499 112301
rect 80010 112296 150499 112298
rect 80010 112240 150438 112296
rect 150494 112240 150499 112296
rect 80010 112238 150499 112240
rect 150433 112235 150499 112238
rect 164693 112298 164759 112301
rect 167494 112298 167500 112300
rect 164693 112296 167500 112298
rect 164693 112240 164698 112296
rect 164754 112240 167500 112296
rect 164693 112238 167500 112240
rect 164693 112235 164759 112238
rect 167494 112236 167500 112238
rect 167564 112236 167570 112300
rect 162025 112162 162091 112165
rect 75134 112160 162091 112162
rect 75134 112104 162030 112160
rect 162086 112104 162091 112160
rect 75134 112102 162091 112104
rect 66069 112099 66135 112102
rect 74993 112099 75059 112102
rect 162025 112099 162091 112102
rect 166993 112162 167059 112165
rect 166993 112160 170292 112162
rect 166993 112104 166998 112160
rect 167054 112104 170292 112160
rect 166993 112102 170292 112104
rect 166993 112099 167059 112102
rect 199694 112100 199700 112164
rect 199764 112100 199770 112164
rect 69422 111964 69428 112028
rect 69492 112026 69498 112028
rect 69492 111966 165354 112026
rect 69492 111964 69498 111966
rect 70158 111828 70164 111892
rect 70228 111890 70234 111892
rect 74993 111890 75059 111893
rect 164693 111890 164759 111893
rect 70228 111830 71146 111890
rect 70228 111828 70234 111830
rect 71086 111754 71146 111830
rect 74993 111888 164759 111890
rect 74993 111832 74998 111888
rect 75054 111832 164698 111888
rect 164754 111832 164759 111888
rect 74993 111830 164759 111832
rect 165294 111890 165354 111966
rect 166901 111890 166967 111893
rect 167310 111890 167316 111892
rect 165294 111888 167316 111890
rect 165294 111832 166906 111888
rect 166962 111832 167316 111888
rect 165294 111830 167316 111832
rect 74993 111827 75059 111830
rect 164693 111827 164759 111830
rect 166901 111827 166967 111830
rect 167310 111828 167316 111830
rect 167380 111828 167386 111892
rect 200062 111828 200068 111892
rect 200132 111890 200138 111892
rect 201861 111890 201927 111893
rect 200132 111888 201927 111890
rect 200132 111832 201866 111888
rect 201922 111832 201927 111888
rect 200132 111830 201927 111832
rect 200132 111828 200138 111830
rect 201861 111827 201927 111830
rect 71086 111694 161490 111754
rect 69841 111618 69907 111621
rect 161430 111618 161490 111694
rect 69841 111616 70380 111618
rect 69841 111560 69846 111616
rect 69902 111560 70380 111616
rect 69841 111558 70380 111560
rect 161430 111558 170292 111618
rect 69841 111555 69907 111558
rect 199694 111420 199700 111484
rect 199764 111420 199770 111484
rect 70158 111284 70164 111348
rect 70228 111346 70234 111348
rect 70228 111286 70410 111346
rect 70228 111284 70234 111286
rect 69054 110876 69060 110940
rect 69124 110938 69130 110940
rect 70350 110938 70410 111286
rect 106038 111148 106044 111212
rect 106108 111210 106114 111212
rect 108941 111210 109007 111213
rect 106108 111208 109007 111210
rect 106108 111152 108946 111208
rect 109002 111152 109007 111208
rect 106108 111150 109007 111152
rect 106108 111148 106114 111150
rect 108941 111147 109007 111150
rect 200062 111148 200068 111212
rect 200132 111210 200138 111212
rect 202045 111210 202111 111213
rect 200132 111208 202111 111210
rect 200132 111152 202050 111208
rect 202106 111152 202111 111208
rect 200132 111150 202111 111152
rect 200132 111148 200138 111150
rect 202045 111147 202111 111150
rect 69124 110908 70410 110938
rect 69124 110878 70380 110908
rect 69124 110876 69130 110878
rect 105670 110876 105676 110940
rect 105740 110876 105746 110940
rect -960 110666 480 110756
rect 169334 110740 169340 110804
rect 169404 110802 169410 110804
rect 169477 110802 169543 110805
rect 169404 110800 170292 110802
rect 169404 110744 169482 110800
rect 169538 110744 170292 110800
rect 169404 110742 170292 110744
rect 169404 110740 169410 110742
rect 169477 110739 169543 110742
rect 199694 110740 199700 110804
rect 199764 110740 199770 110804
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 200062 110468 200068 110532
rect 200132 110530 200138 110532
rect 200389 110530 200455 110533
rect 200132 110528 200455 110530
rect 200132 110472 200394 110528
rect 200450 110472 200455 110528
rect 200132 110470 200455 110472
rect 200132 110468 200138 110470
rect 200389 110467 200455 110470
rect 106038 110332 106044 110396
rect 106108 110394 106114 110396
rect 108941 110394 109007 110397
rect 106108 110392 109007 110394
rect 106108 110336 108946 110392
rect 109002 110336 109007 110392
rect 106108 110334 109007 110336
rect 106108 110332 106114 110334
rect 108941 110331 109007 110334
rect 105670 110196 105676 110260
rect 105740 110196 105746 110260
rect 166993 110258 167059 110261
rect 166993 110256 170292 110258
rect 166993 110200 166998 110256
rect 167054 110200 170292 110256
rect 166993 110198 170292 110200
rect 166993 110195 167059 110198
rect 199694 110060 199700 110124
rect 199764 110060 199770 110124
rect 70301 109986 70367 109989
rect 70301 109984 70410 109986
rect 70301 109928 70306 109984
rect 70362 109928 70410 109984
rect 70301 109923 70410 109928
rect 70350 109548 70410 109923
rect 106038 109788 106044 109852
rect 106108 109850 106114 109852
rect 108573 109850 108639 109853
rect 106108 109848 108639 109850
rect 106108 109792 108578 109848
rect 108634 109792 108639 109848
rect 106108 109790 108639 109792
rect 106108 109788 106114 109790
rect 108573 109787 108639 109790
rect 200062 109788 200068 109852
rect 200132 109850 200138 109852
rect 201861 109850 201927 109853
rect 200132 109848 201927 109850
rect 200132 109792 201866 109848
rect 201922 109792 201927 109848
rect 200132 109790 201927 109792
rect 200132 109788 200138 109790
rect 201861 109787 201927 109790
rect 105670 109516 105676 109580
rect 105740 109516 105746 109580
rect 167085 109578 167151 109581
rect 169385 109578 169451 109581
rect 167085 109576 170292 109578
rect 167085 109520 167090 109576
rect 167146 109520 169390 109576
rect 169446 109520 170292 109576
rect 167085 109518 170292 109520
rect 167085 109515 167151 109518
rect 169385 109515 169451 109518
rect 199694 109380 199700 109444
rect 199764 109380 199770 109444
rect 200062 109108 200068 109172
rect 200132 109170 200138 109172
rect 202781 109170 202847 109173
rect 200132 109168 202847 109170
rect 200132 109112 202786 109168
rect 202842 109112 202847 109168
rect 200132 109110 202847 109112
rect 200132 109108 200138 109110
rect 202781 109107 202847 109110
rect 106038 108972 106044 109036
rect 106108 109034 106114 109036
rect 107653 109034 107719 109037
rect 106108 109032 107719 109034
rect 106108 108976 107658 109032
rect 107714 108976 107719 109032
rect 106108 108974 107719 108976
rect 106108 108972 106114 108974
rect 107653 108971 107719 108974
rect 70342 108836 70348 108900
rect 70412 108836 70418 108900
rect 105670 108836 105676 108900
rect 105740 108836 105746 108900
rect 168925 108898 168991 108901
rect 169886 108898 169892 108900
rect 168925 108896 169892 108898
rect 168925 108840 168930 108896
rect 168986 108840 169892 108896
rect 168925 108838 169892 108840
rect 168925 108835 168991 108838
rect 169886 108836 169892 108838
rect 169956 108898 169962 108900
rect 169956 108838 170292 108898
rect 169956 108836 169962 108838
rect 70209 108626 70275 108629
rect 70209 108624 70410 108626
rect 70209 108568 70214 108624
rect 70270 108568 70410 108624
rect 70209 108566 70410 108568
rect 70209 108563 70275 108566
rect 70350 108188 70410 108566
rect 106038 108428 106044 108492
rect 106108 108490 106114 108492
rect 106365 108490 106431 108493
rect 108021 108490 108087 108493
rect 106108 108488 108087 108490
rect 106108 108432 106370 108488
rect 106426 108432 108026 108488
rect 108082 108432 108087 108488
rect 106108 108430 108087 108432
rect 106108 108428 106114 108430
rect 106365 108427 106431 108430
rect 108021 108427 108087 108430
rect 200062 108428 200068 108492
rect 200132 108490 200138 108492
rect 200297 108490 200363 108493
rect 200132 108488 200363 108490
rect 200132 108432 200302 108488
rect 200358 108432 200363 108488
rect 200132 108430 200363 108432
rect 200132 108428 200138 108430
rect 200297 108427 200363 108430
rect 105670 108156 105676 108220
rect 105740 108156 105746 108220
rect 199694 108156 199700 108220
rect 199764 108156 199770 108220
rect 68829 107538 68895 107541
rect 166993 107538 167059 107541
rect 68829 107536 70380 107538
rect 68829 107480 68834 107536
rect 68890 107480 70380 107536
rect 68829 107478 70380 107480
rect 166993 107536 170292 107538
rect 166993 107480 166998 107536
rect 167054 107480 170292 107536
rect 166993 107478 170292 107480
rect 68829 107475 68895 107478
rect 166993 107475 167059 107478
rect 105670 107340 105676 107404
rect 105740 107340 105746 107404
rect 199694 107340 199700 107404
rect 199764 107340 199770 107404
rect 106038 107068 106044 107132
rect 106108 107130 106114 107132
rect 108941 107130 109007 107133
rect 106108 107128 109007 107130
rect 106108 107072 108946 107128
rect 109002 107072 109007 107128
rect 106108 107070 109007 107072
rect 106108 107068 106114 107070
rect 108941 107067 109007 107070
rect 200062 107068 200068 107132
rect 200132 107130 200138 107132
rect 202781 107130 202847 107133
rect 200132 107128 202847 107130
rect 200132 107072 202786 107128
rect 202842 107072 202847 107128
rect 200132 107070 202847 107072
rect 200132 107068 200138 107070
rect 202781 107067 202847 107070
rect 68553 106858 68619 106861
rect 68553 106856 70380 106858
rect 68553 106800 68558 106856
rect 68614 106800 70380 106856
rect 68553 106798 70380 106800
rect 68553 106795 68619 106798
rect 105670 106660 105676 106724
rect 105740 106660 105746 106724
rect 166993 106722 167059 106725
rect 166993 106720 170292 106722
rect 166993 106664 166998 106720
rect 167054 106664 170292 106720
rect 166993 106662 170292 106664
rect 166993 106659 167059 106662
rect 199694 106660 199700 106724
rect 199764 106660 199770 106724
rect 106038 106388 106044 106452
rect 106108 106450 106114 106452
rect 108941 106450 109007 106453
rect 106108 106448 109007 106450
rect 106108 106392 108946 106448
rect 109002 106392 109007 106448
rect 106108 106390 109007 106392
rect 106108 106388 106114 106390
rect 108941 106387 109007 106390
rect 200062 106388 200068 106452
rect 200132 106450 200138 106452
rect 202229 106450 202295 106453
rect 200132 106448 202295 106450
rect 200132 106392 202234 106448
rect 202290 106392 202295 106448
rect 200132 106390 202295 106392
rect 200132 106388 200138 106390
rect 202229 106387 202295 106390
rect 169109 106178 169175 106181
rect 169845 106178 169911 106181
rect 169109 106176 170292 106178
rect 169109 106120 169114 106176
rect 169170 106120 169850 106176
rect 169906 106120 170292 106176
rect 169109 106118 170292 106120
rect 169109 106115 169175 106118
rect 169845 106115 169911 106118
rect 69105 106042 69171 106045
rect 69105 106040 70380 106042
rect 69105 105984 69110 106040
rect 69166 105984 70380 106040
rect 69105 105982 70380 105984
rect 69105 105979 69171 105982
rect 105670 105980 105676 106044
rect 105740 105980 105746 106044
rect 199510 105980 199516 106044
rect 199580 105980 199586 106044
rect 106038 105708 106044 105772
rect 106108 105770 106114 105772
rect 108941 105770 109007 105773
rect 106108 105768 109007 105770
rect 106108 105712 108946 105768
rect 109002 105712 109007 105768
rect 106108 105710 109007 105712
rect 106108 105708 106114 105710
rect 108941 105707 109007 105710
rect 200062 105708 200068 105772
rect 200132 105770 200138 105772
rect 201585 105770 201651 105773
rect 200132 105768 201651 105770
rect 200132 105712 201590 105768
rect 201646 105712 201651 105768
rect 200132 105710 201651 105712
rect 200132 105708 200138 105710
rect 201585 105707 201651 105710
rect 67541 105498 67607 105501
rect 167913 105498 167979 105501
rect 67541 105496 70380 105498
rect 67541 105440 67546 105496
rect 67602 105440 70380 105496
rect 67541 105438 70380 105440
rect 167913 105496 170292 105498
rect 167913 105440 167918 105496
rect 167974 105440 170292 105496
rect 167913 105438 170292 105440
rect 67541 105435 67607 105438
rect 167913 105435 167979 105438
rect 199694 105436 199700 105500
rect 199764 105436 199770 105500
rect 200062 105028 200068 105092
rect 200132 105090 200138 105092
rect 201769 105090 201835 105093
rect 200132 105088 201835 105090
rect 200132 105032 201774 105088
rect 201830 105032 201835 105088
rect 200132 105030 201835 105032
rect 200132 105028 200138 105030
rect 201769 105027 201835 105030
rect 67633 104818 67699 104821
rect 67633 104816 70380 104818
rect 67633 104760 67638 104816
rect 67694 104760 70380 104816
rect 67633 104758 70380 104760
rect 67633 104755 67699 104758
rect 105670 104756 105676 104820
rect 105740 104756 105746 104820
rect 106038 104756 106044 104820
rect 106108 104818 106114 104820
rect 106457 104818 106523 104821
rect 108021 104818 108087 104821
rect 106108 104816 108087 104818
rect 106108 104760 106462 104816
rect 106518 104760 108026 104816
rect 108082 104760 108087 104816
rect 106108 104758 108087 104760
rect 106108 104756 106114 104758
rect 106457 104755 106523 104758
rect 108021 104755 108087 104758
rect 169017 104818 169083 104821
rect 169017 104816 170292 104818
rect 169017 104760 169022 104816
rect 169078 104760 170292 104816
rect 169017 104758 170292 104760
rect 169017 104755 169083 104758
rect 199510 104620 199516 104684
rect 199580 104620 199586 104684
rect 106038 104348 106044 104412
rect 106108 104410 106114 104412
rect 108205 104410 108271 104413
rect 200113 104412 200179 104413
rect 106108 104408 108271 104410
rect 106108 104352 108210 104408
rect 108266 104352 108271 104408
rect 106108 104350 108271 104352
rect 106108 104348 106114 104350
rect 108205 104347 108271 104350
rect 200062 104348 200068 104412
rect 200132 104410 200179 104412
rect 200132 104408 200224 104410
rect 200174 104352 200224 104408
rect 200132 104350 200224 104352
rect 200132 104348 200179 104350
rect 200113 104347 200179 104348
rect 66989 104138 67055 104141
rect 66989 104136 70380 104138
rect 66989 104080 66994 104136
rect 67050 104080 70380 104136
rect 66989 104078 70380 104080
rect 66989 104075 67055 104078
rect 105670 104076 105676 104140
rect 105740 104076 105746 104140
rect 169201 104138 169267 104141
rect 169201 104136 170292 104138
rect 169201 104080 169206 104136
rect 169262 104080 170292 104136
rect 169201 104078 170292 104080
rect 169201 104075 169267 104078
rect 199694 104076 199700 104140
rect 199764 104076 199770 104140
rect 200062 103668 200068 103732
rect 200132 103730 200138 103732
rect 201861 103730 201927 103733
rect 200132 103728 201927 103730
rect 200132 103672 201866 103728
rect 201922 103672 201927 103728
rect 200132 103670 201927 103672
rect 200132 103668 200138 103670
rect 201861 103667 201927 103670
rect 166993 103458 167059 103461
rect 166993 103456 170292 103458
rect 166993 103400 166998 103456
rect 167054 103400 170292 103456
rect 166993 103398 170292 103400
rect 166993 103395 167059 103398
rect 105670 103260 105676 103324
rect 105740 103260 105746 103324
rect 106038 102988 106044 103052
rect 106108 103050 106114 103052
rect 108941 103050 109007 103053
rect 106108 103048 109007 103050
rect 106108 102992 108946 103048
rect 109002 102992 109007 103048
rect 106108 102990 109007 102992
rect 106108 102988 106114 102990
rect 108941 102987 109007 102990
rect 200062 102988 200068 103052
rect 200132 103050 200138 103052
rect 201677 103050 201743 103053
rect 200132 103048 201743 103050
rect 200132 102992 201682 103048
rect 201738 102992 201743 103048
rect 200132 102990 201743 102992
rect 200132 102988 200138 102990
rect 201677 102987 201743 102990
rect 67633 102778 67699 102781
rect 67633 102776 70380 102778
rect 67633 102720 67638 102776
rect 67694 102720 70380 102776
rect 67633 102718 70380 102720
rect 67633 102715 67699 102718
rect 199694 102716 199700 102780
rect 199764 102716 199770 102780
rect 105670 102580 105676 102644
rect 105740 102580 105746 102644
rect 106038 102308 106044 102372
rect 106108 102370 106114 102372
rect 106457 102370 106523 102373
rect 108205 102370 108271 102373
rect 106108 102368 108271 102370
rect 106108 102312 106462 102368
rect 106518 102312 108210 102368
rect 108266 102312 108271 102368
rect 106108 102310 108271 102312
rect 106108 102308 106114 102310
rect 106457 102307 106523 102310
rect 108205 102307 108271 102310
rect 67214 102036 67220 102100
rect 67284 102098 67290 102100
rect 166993 102098 167059 102101
rect 67284 102038 70380 102098
rect 166993 102096 170292 102098
rect 166993 102040 166998 102096
rect 167054 102040 170292 102096
rect 166993 102038 170292 102040
rect 67284 102036 67290 102038
rect 166993 102035 167059 102038
rect 105670 101900 105676 101964
rect 105740 101900 105746 101964
rect 199694 101900 199700 101964
rect 199764 101900 199770 101964
rect 106038 101628 106044 101692
rect 106108 101690 106114 101692
rect 108941 101690 109007 101693
rect 106108 101688 109007 101690
rect 106108 101632 108946 101688
rect 109002 101632 109007 101688
rect 106108 101630 109007 101632
rect 106108 101628 106114 101630
rect 108941 101627 109007 101630
rect 200062 101628 200068 101692
rect 200132 101690 200138 101692
rect 201861 101690 201927 101693
rect 200132 101688 201927 101690
rect 200132 101632 201866 101688
rect 201922 101632 201927 101688
rect 200132 101630 201927 101632
rect 200132 101628 200138 101630
rect 201861 101627 201927 101630
rect 67265 101418 67331 101421
rect 67265 101416 70380 101418
rect 67265 101360 67270 101416
rect 67326 101360 70380 101416
rect 67265 101358 70380 101360
rect 67265 101355 67331 101358
rect 105670 101220 105676 101284
rect 105740 101220 105746 101284
rect 167494 101220 167500 101284
rect 167564 101282 167570 101284
rect 169518 101282 169524 101284
rect 167564 101222 169524 101282
rect 167564 101220 167570 101222
rect 169518 101220 169524 101222
rect 169588 101282 169594 101284
rect 169588 101222 170292 101282
rect 169588 101220 169594 101222
rect 199694 101220 199700 101284
rect 199764 101220 199770 101284
rect 106038 100948 106044 101012
rect 106108 101010 106114 101012
rect 108757 101010 108823 101013
rect 106108 101008 108823 101010
rect 106108 100952 108762 101008
rect 108818 100952 108823 101008
rect 106108 100950 108823 100952
rect 106108 100948 106114 100950
rect 108757 100947 108823 100950
rect 200062 100948 200068 101012
rect 200132 101010 200138 101012
rect 201534 101010 201540 101012
rect 200132 100950 201540 101010
rect 200132 100948 200138 100950
rect 201534 100948 201540 100950
rect 201604 100948 201610 101012
rect 67633 100738 67699 100741
rect 167453 100738 167519 100741
rect 169017 100738 169083 100741
rect 67633 100736 70380 100738
rect 67633 100680 67638 100736
rect 67694 100680 70380 100736
rect 67633 100678 70380 100680
rect 167453 100736 170292 100738
rect 167453 100680 167458 100736
rect 167514 100680 169022 100736
rect 169078 100680 170292 100736
rect 167453 100678 170292 100680
rect 67633 100675 67699 100678
rect 167453 100675 167519 100678
rect 169017 100675 169083 100678
rect 105670 100540 105676 100604
rect 105740 100540 105746 100604
rect 199694 100540 199700 100604
rect 199764 100540 199770 100604
rect 106038 100268 106044 100332
rect 106108 100330 106114 100332
rect 108941 100330 109007 100333
rect 106108 100328 109007 100330
rect 106108 100272 108946 100328
rect 109002 100272 109007 100328
rect 106108 100270 109007 100272
rect 106108 100268 106114 100270
rect 108941 100267 109007 100270
rect 200062 100268 200068 100332
rect 200132 100330 200138 100332
rect 201585 100330 201651 100333
rect 200132 100328 201651 100330
rect 200132 100272 201590 100328
rect 201646 100272 201651 100328
rect 200132 100270 201651 100272
rect 200132 100268 200138 100270
rect 201585 100267 201651 100270
rect 68277 100058 68343 100061
rect 167085 100058 167151 100061
rect 169477 100058 169543 100061
rect 68277 100056 70380 100058
rect 68277 100000 68282 100056
rect 68338 100000 70380 100056
rect 68277 99998 70380 100000
rect 167085 100056 170292 100058
rect 167085 100000 167090 100056
rect 167146 100000 169482 100056
rect 169538 100000 170292 100056
rect 167085 99998 170292 100000
rect 68277 99995 68343 99998
rect 167085 99995 167151 99998
rect 169477 99995 169543 99998
rect 105670 99860 105676 99924
rect 105740 99860 105746 99924
rect 199694 99860 199700 99924
rect 199764 99860 199770 99924
rect 106038 99588 106044 99652
rect 106108 99650 106114 99652
rect 108757 99650 108823 99653
rect 106108 99648 108823 99650
rect 106108 99592 108762 99648
rect 108818 99592 108823 99648
rect 106108 99590 108823 99592
rect 106108 99588 106114 99590
rect 108757 99587 108823 99590
rect 200062 99588 200068 99652
rect 200132 99650 200138 99652
rect 202781 99650 202847 99653
rect 200132 99648 202847 99650
rect 200132 99592 202786 99648
rect 202842 99592 202847 99648
rect 200132 99590 202847 99592
rect 200132 99588 200138 99590
rect 202781 99587 202847 99590
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 69565 99378 69631 99381
rect 69565 99376 70380 99378
rect 69565 99320 69570 99376
rect 69626 99320 70380 99376
rect 583520 99364 584960 99454
rect 69565 99318 70380 99320
rect 69565 99315 69631 99318
rect 105670 99180 105676 99244
rect 105740 99180 105746 99244
rect 106038 98908 106044 98972
rect 106108 98970 106114 98972
rect 107653 98970 107719 98973
rect 170070 98970 170076 98972
rect 106108 98968 107719 98970
rect 106108 98912 107658 98968
rect 107714 98912 107719 98968
rect 106108 98910 107719 98912
rect 106108 98908 106114 98910
rect 107653 98907 107719 98910
rect 161430 98910 170076 98970
rect 67633 98698 67699 98701
rect 67633 98696 70380 98698
rect 67633 98640 67638 98696
rect 67694 98640 70380 98696
rect 67633 98638 70380 98640
rect 67633 98635 67699 98638
rect 145557 98018 145623 98021
rect 161430 98018 161490 98910
rect 170070 98908 170076 98910
rect 170140 98970 170146 98972
rect 170262 98970 170322 99212
rect 199694 99180 199700 99244
rect 199764 99180 199770 99244
rect 170140 98910 170322 98970
rect 170140 98908 170146 98910
rect 200062 98908 200068 98972
rect 200132 98970 200138 98972
rect 201585 98970 201651 98973
rect 200132 98968 201651 98970
rect 200132 98912 201590 98968
rect 201646 98912 201651 98968
rect 200132 98910 201651 98912
rect 200132 98908 200138 98910
rect 201585 98907 201651 98910
rect 167545 98698 167611 98701
rect 169109 98698 169175 98701
rect 167545 98696 170292 98698
rect 167545 98640 167550 98696
rect 167606 98640 169114 98696
rect 169170 98640 170292 98696
rect 167545 98638 170292 98640
rect 167545 98635 167611 98638
rect 169109 98635 169175 98638
rect 199694 98500 199700 98564
rect 199764 98500 199770 98564
rect 200113 98292 200179 98293
rect 200062 98228 200068 98292
rect 200132 98290 200179 98292
rect 200132 98288 200224 98290
rect 200174 98232 200224 98288
rect 200132 98230 200224 98232
rect 200132 98228 200179 98230
rect 200113 98227 200179 98228
rect 145557 98016 161490 98018
rect 145557 97960 145562 98016
rect 145618 97960 161490 98016
rect 145557 97958 161490 97960
rect 145557 97955 145623 97958
rect 67633 97882 67699 97885
rect 67633 97880 70380 97882
rect 67633 97824 67638 97880
rect 67694 97824 70380 97880
rect 67633 97822 70380 97824
rect 67633 97819 67699 97822
rect 105670 97820 105676 97884
rect 105740 97820 105746 97884
rect 106038 97820 106044 97884
rect 106108 97882 106114 97884
rect 106549 97882 106615 97885
rect 107745 97882 107811 97885
rect 106108 97880 107811 97882
rect 106108 97824 106554 97880
rect 106610 97824 107750 97880
rect 107806 97824 107811 97880
rect 106108 97822 107811 97824
rect 106108 97820 106114 97822
rect 106549 97819 106615 97822
rect 107745 97819 107811 97822
rect 167177 97882 167243 97885
rect 168925 97882 168991 97885
rect 167177 97880 170292 97882
rect 167177 97824 167182 97880
rect 167238 97824 168930 97880
rect 168986 97824 170292 97880
rect 167177 97822 170292 97824
rect 167177 97819 167243 97822
rect 168925 97819 168991 97822
rect -960 97610 480 97700
rect 3601 97610 3667 97613
rect -960 97608 3667 97610
rect -960 97552 3606 97608
rect 3662 97552 3667 97608
rect -960 97550 3667 97552
rect -960 97460 480 97550
rect 3601 97547 3667 97550
rect 106038 97548 106044 97612
rect 106108 97610 106114 97612
rect 107653 97610 107719 97613
rect 106108 97608 107719 97610
rect 106108 97552 107658 97608
rect 107714 97552 107719 97608
rect 106108 97550 107719 97552
rect 106108 97548 106114 97550
rect 107653 97547 107719 97550
rect 200062 97548 200068 97612
rect 200132 97610 200138 97612
rect 201953 97610 202019 97613
rect 200132 97608 202019 97610
rect 200132 97552 201958 97608
rect 202014 97552 202019 97608
rect 200132 97550 202019 97552
rect 200132 97548 200138 97550
rect 201953 97547 202019 97550
rect 69657 97338 69723 97341
rect 69657 97336 70380 97338
rect 69657 97280 69662 97336
rect 69718 97280 70380 97336
rect 69657 97278 70380 97280
rect 69657 97275 69723 97278
rect 105486 97276 105492 97340
rect 105556 97276 105562 97340
rect 199694 97276 199700 97340
rect 199764 97276 199770 97340
rect 200062 96868 200068 96932
rect 200132 96868 200138 96932
rect 105670 96596 105676 96660
rect 105740 96596 105746 96660
rect 199694 96596 199700 96660
rect 199764 96596 199770 96660
rect 106038 96460 106044 96524
rect 106108 96522 106114 96524
rect 107745 96522 107811 96525
rect 106108 96520 107811 96522
rect 106108 96464 107750 96520
rect 107806 96464 107811 96520
rect 106108 96462 107811 96464
rect 106108 96460 106114 96462
rect 107745 96459 107811 96462
rect 162669 96522 162735 96525
rect 167494 96522 167500 96524
rect 162669 96520 167500 96522
rect 162669 96464 162674 96520
rect 162730 96464 167500 96520
rect 162669 96462 167500 96464
rect 162669 96459 162735 96462
rect 167494 96460 167500 96462
rect 167564 96522 167570 96524
rect 200070 96522 200130 96868
rect 202137 96522 202203 96525
rect 167564 96462 170292 96522
rect 200070 96520 202203 96522
rect 200070 96464 202142 96520
rect 202198 96464 202203 96520
rect 200070 96462 202203 96464
rect 167564 96460 167570 96462
rect 202137 96459 202203 96462
rect 106038 96188 106044 96252
rect 106108 96250 106114 96252
rect 107653 96250 107719 96253
rect 106108 96248 107719 96250
rect 106108 96192 107658 96248
rect 107714 96192 107719 96248
rect 106108 96190 107719 96192
rect 106108 96188 106114 96190
rect 107653 96187 107719 96190
rect 200062 96188 200068 96252
rect 200132 96250 200138 96252
rect 202413 96250 202479 96253
rect 200132 96248 202479 96250
rect 200132 96192 202418 96248
rect 202474 96192 202479 96248
rect 200132 96190 202479 96192
rect 200132 96188 200138 96190
rect 202413 96187 202479 96190
rect 67633 95978 67699 95981
rect 67633 95976 70380 95978
rect 67633 95920 67638 95976
rect 67694 95920 70380 95976
rect 67633 95918 70380 95920
rect 67633 95915 67699 95918
rect 105670 95916 105676 95980
rect 105740 95916 105746 95980
rect 199694 95916 199700 95980
rect 199764 95916 199770 95980
rect 167310 95780 167316 95844
rect 167380 95842 167386 95844
rect 167380 95782 170292 95842
rect 167380 95780 167386 95782
rect 106038 95508 106044 95572
rect 106108 95570 106114 95572
rect 107837 95570 107903 95573
rect 106108 95568 107903 95570
rect 106108 95512 107842 95568
rect 107898 95512 107903 95568
rect 106108 95510 107903 95512
rect 106108 95508 106114 95510
rect 107837 95507 107903 95510
rect 200062 95508 200068 95572
rect 200132 95570 200138 95572
rect 200205 95570 200271 95573
rect 201401 95570 201467 95573
rect 200132 95568 201467 95570
rect 200132 95512 200210 95568
rect 200266 95512 201406 95568
rect 201462 95512 201467 95568
rect 200132 95510 201467 95512
rect 200132 95508 200138 95510
rect 200205 95507 200271 95510
rect 201401 95507 201467 95510
rect 69197 95298 69263 95301
rect 119981 95300 120047 95301
rect 69197 95296 70380 95298
rect 69197 95240 69202 95296
rect 69258 95240 70380 95296
rect 69197 95238 70380 95240
rect 69197 95235 69263 95238
rect 105670 95236 105676 95300
rect 105740 95236 105746 95300
rect 119981 95296 120028 95300
rect 120092 95298 120098 95300
rect 168833 95298 168899 95301
rect 119981 95240 119986 95296
rect 119981 95236 120028 95240
rect 120092 95238 120138 95298
rect 168833 95296 170292 95298
rect 168833 95240 168838 95296
rect 168894 95240 170292 95296
rect 168833 95238 170292 95240
rect 120092 95236 120098 95238
rect 119981 95235 120047 95236
rect 168833 95235 168899 95238
rect 199694 95236 199700 95300
rect 199764 95236 199770 95300
rect 106038 94828 106044 94892
rect 106108 94890 106114 94892
rect 107653 94890 107719 94893
rect 106108 94888 107719 94890
rect 106108 94832 107658 94888
rect 107714 94832 107719 94888
rect 106108 94830 107719 94832
rect 106108 94828 106114 94830
rect 107653 94827 107719 94830
rect 200062 94828 200068 94892
rect 200132 94890 200138 94892
rect 200205 94890 200271 94893
rect 200132 94888 200271 94890
rect 200132 94832 200210 94888
rect 200266 94832 200271 94888
rect 200132 94830 200271 94832
rect 200132 94828 200138 94830
rect 200205 94827 200271 94830
rect 68921 94618 68987 94621
rect 166993 94618 167059 94621
rect 68921 94616 70380 94618
rect 68921 94560 68926 94616
rect 68982 94560 70380 94616
rect 68921 94558 70380 94560
rect 166993 94616 170292 94618
rect 166993 94560 166998 94616
rect 167054 94560 170292 94616
rect 166993 94558 170292 94560
rect 68921 94555 68987 94558
rect 166993 94555 167059 94558
rect 199694 94556 199700 94620
rect 199764 94556 199770 94620
rect 105670 94420 105676 94484
rect 105740 94420 105746 94484
rect 106038 94148 106044 94212
rect 106108 94210 106114 94212
rect 107653 94210 107719 94213
rect 106108 94208 107719 94210
rect 106108 94152 107658 94208
rect 107714 94152 107719 94208
rect 106108 94150 107719 94152
rect 106108 94148 106114 94150
rect 107653 94147 107719 94150
rect 200062 94148 200068 94212
rect 200132 94210 200138 94212
rect 202781 94210 202847 94213
rect 200132 94208 202847 94210
rect 200132 94152 202786 94208
rect 202842 94152 202847 94208
rect 200132 94150 202847 94152
rect 200132 94148 200138 94150
rect 202781 94147 202847 94150
rect 69473 93938 69539 93941
rect 69473 93936 70380 93938
rect 69473 93880 69478 93936
rect 69534 93880 70380 93936
rect 69473 93878 70380 93880
rect 69473 93875 69539 93878
rect 105486 93876 105492 93940
rect 105556 93876 105562 93940
rect 167729 93938 167795 93941
rect 167729 93936 170292 93938
rect 167729 93880 167734 93936
rect 167790 93880 170292 93936
rect 167729 93878 170292 93880
rect 167729 93875 167795 93878
rect 199694 93876 199700 93940
rect 199764 93876 199770 93940
rect 106038 93468 106044 93532
rect 106108 93530 106114 93532
rect 107653 93530 107719 93533
rect 106108 93528 107719 93530
rect 106108 93472 107658 93528
rect 107714 93472 107719 93528
rect 106108 93470 107719 93472
rect 106108 93468 106114 93470
rect 107653 93467 107719 93470
rect 67633 93258 67699 93261
rect 67633 93256 70380 93258
rect 67633 93200 67638 93256
rect 67694 93200 70380 93256
rect 67633 93198 70380 93200
rect 67633 93195 67699 93198
rect 105670 93196 105676 93260
rect 105740 93196 105746 93260
rect 166901 93258 166967 93261
rect 166901 93256 170292 93258
rect 166901 93200 166906 93256
rect 166962 93200 170292 93256
rect 166901 93198 170292 93200
rect 166901 93195 166967 93198
rect 199694 93060 199700 93124
rect 199764 93060 199770 93124
rect 106038 92788 106044 92852
rect 106108 92850 106114 92852
rect 107745 92850 107811 92853
rect 106108 92848 107811 92850
rect 106108 92792 107750 92848
rect 107806 92792 107811 92848
rect 106108 92790 107811 92792
rect 106108 92788 106114 92790
rect 107745 92787 107811 92790
rect 200062 92788 200068 92852
rect 200132 92850 200138 92852
rect 200297 92850 200363 92853
rect 200132 92848 200363 92850
rect 200132 92792 200302 92848
rect 200358 92792 200363 92848
rect 200132 92790 200363 92792
rect 200132 92788 200138 92790
rect 200297 92787 200363 92790
rect 69422 92516 69428 92580
rect 69492 92578 69498 92580
rect 69492 92518 70380 92578
rect 69492 92516 69498 92518
rect 105670 92516 105676 92580
rect 105740 92516 105746 92580
rect 167269 92578 167335 92581
rect 167913 92578 167979 92581
rect 167269 92576 170292 92578
rect 167269 92520 167274 92576
rect 167330 92520 167918 92576
rect 167974 92520 170292 92576
rect 167269 92518 170292 92520
rect 167269 92515 167335 92518
rect 167913 92515 167979 92518
rect 200062 92108 200068 92172
rect 200132 92170 200138 92172
rect 202045 92170 202111 92173
rect 200132 92168 202111 92170
rect 200132 92112 202050 92168
rect 202106 92112 202111 92168
rect 200132 92110 202111 92112
rect 200132 92108 200138 92110
rect 202045 92107 202111 92110
rect 68093 91898 68159 91901
rect 68093 91896 70380 91898
rect 68093 91840 68098 91896
rect 68154 91840 70380 91896
rect 68093 91838 70380 91840
rect 68093 91835 68159 91838
rect 199694 91836 199700 91900
rect 199764 91836 199770 91900
rect 106038 91428 106044 91492
rect 106108 91490 106114 91492
rect 107745 91490 107811 91493
rect 106108 91488 107811 91490
rect 106108 91432 107750 91488
rect 107806 91432 107811 91488
rect 106108 91430 107811 91432
rect 106108 91428 106114 91430
rect 107745 91427 107811 91430
rect 200062 91428 200068 91492
rect 200132 91490 200138 91492
rect 201718 91490 201724 91492
rect 200132 91430 201724 91490
rect 200132 91428 200138 91430
rect 201718 91428 201724 91430
rect 201788 91428 201794 91492
rect 67633 91218 67699 91221
rect 67633 91216 70380 91218
rect 67633 91160 67638 91216
rect 67694 91160 70380 91216
rect 67633 91158 70380 91160
rect 67633 91155 67699 91158
rect 105670 91156 105676 91220
rect 105740 91156 105746 91220
rect 167729 91218 167795 91221
rect 167729 91216 170292 91218
rect 167729 91160 167734 91216
rect 167790 91160 170292 91216
rect 167729 91158 170292 91160
rect 167729 91155 167795 91158
rect 199694 91156 199700 91220
rect 199764 91156 199770 91220
rect 106038 90748 106044 90812
rect 106108 90810 106114 90812
rect 108021 90810 108087 90813
rect 106108 90808 108087 90810
rect 106108 90752 108026 90808
rect 108082 90752 108087 90808
rect 106108 90750 108087 90752
rect 106108 90748 106114 90750
rect 108021 90747 108087 90750
rect 200062 90748 200068 90812
rect 200132 90810 200138 90812
rect 201769 90810 201835 90813
rect 200132 90808 201835 90810
rect 200132 90752 201774 90808
rect 201830 90752 201835 90808
rect 200132 90750 201835 90752
rect 200132 90748 200138 90750
rect 201769 90747 201835 90750
rect 69381 90538 69447 90541
rect 69381 90536 70380 90538
rect 69381 90480 69386 90536
rect 69442 90480 70380 90536
rect 69381 90478 70380 90480
rect 69381 90475 69447 90478
rect 105670 90476 105676 90540
rect 105740 90476 105746 90540
rect 167637 90538 167703 90541
rect 167637 90536 170292 90538
rect 167637 90480 167642 90536
rect 167698 90480 170292 90536
rect 167637 90478 170292 90480
rect 167637 90475 167703 90478
rect 199694 90476 199700 90540
rect 199764 90476 199770 90540
rect 106038 90068 106044 90132
rect 106108 90130 106114 90132
rect 107653 90130 107719 90133
rect 106108 90128 107719 90130
rect 106108 90072 107658 90128
rect 107714 90072 107719 90128
rect 106108 90070 107719 90072
rect 106108 90068 106114 90070
rect 107653 90067 107719 90070
rect 200062 90068 200068 90132
rect 200132 90130 200138 90132
rect 201769 90130 201835 90133
rect 200132 90128 201835 90130
rect 200132 90072 201774 90128
rect 201830 90072 201835 90128
rect 200132 90070 201835 90072
rect 200132 90068 200138 90070
rect 201769 90067 201835 90070
rect 105670 89796 105676 89860
rect 105740 89796 105746 89860
rect 166993 89858 167059 89861
rect 166993 89856 170292 89858
rect 166993 89800 166998 89856
rect 167054 89800 170292 89856
rect 166993 89798 170292 89800
rect 166993 89795 167059 89798
rect 199694 89796 199700 89860
rect 199764 89796 199770 89860
rect 106038 89388 106044 89452
rect 106108 89450 106114 89452
rect 108665 89450 108731 89453
rect 106108 89448 108731 89450
rect 106108 89392 108670 89448
rect 108726 89392 108731 89448
rect 106108 89390 108731 89392
rect 106108 89388 106114 89390
rect 108665 89387 108731 89390
rect 200062 89388 200068 89452
rect 200132 89450 200138 89452
rect 202137 89450 202203 89453
rect 200132 89448 202203 89450
rect 200132 89392 202142 89448
rect 202198 89392 202203 89448
rect 200132 89390 202203 89392
rect 200132 89388 200138 89390
rect 202137 89387 202203 89390
rect 105670 89116 105676 89180
rect 105740 89116 105746 89180
rect 199694 89116 199700 89180
rect 199764 89116 199770 89180
rect 68553 89042 68619 89045
rect 69013 89042 69079 89045
rect 166993 89042 167059 89045
rect 68553 89040 70380 89042
rect 68553 88984 68558 89040
rect 68614 88984 69018 89040
rect 69074 88984 70380 89040
rect 68553 88982 70380 88984
rect 166993 89040 170292 89042
rect 166993 88984 166998 89040
rect 167054 88984 170292 89040
rect 166993 88982 170292 88984
rect 68553 88979 68619 88982
rect 69013 88979 69079 88982
rect 166993 88979 167059 88982
rect 106038 88708 106044 88772
rect 106108 88770 106114 88772
rect 108573 88770 108639 88773
rect 106108 88768 108639 88770
rect 106108 88712 108578 88768
rect 108634 88712 108639 88768
rect 106108 88710 108639 88712
rect 106108 88708 106114 88710
rect 108573 88707 108639 88710
rect 200062 88708 200068 88772
rect 200132 88770 200138 88772
rect 202505 88770 202571 88773
rect 200132 88768 202571 88770
rect 200132 88712 202510 88768
rect 202566 88712 202571 88768
rect 200132 88710 202571 88712
rect 200132 88708 200138 88710
rect 202505 88707 202571 88710
rect 68461 88498 68527 88501
rect 68461 88496 70380 88498
rect 68461 88440 68466 88496
rect 68522 88440 70380 88496
rect 68461 88438 70380 88440
rect 68461 88435 68527 88438
rect 105670 88436 105676 88500
rect 105740 88436 105746 88500
rect 167177 88498 167243 88501
rect 169753 88498 169819 88501
rect 167177 88496 170292 88498
rect 167177 88440 167182 88496
rect 167238 88440 169758 88496
rect 169814 88440 170292 88496
rect 167177 88438 170292 88440
rect 167177 88435 167243 88438
rect 169753 88435 169819 88438
rect 199694 88436 199700 88500
rect 199764 88436 199770 88500
rect 106038 88028 106044 88092
rect 106108 88090 106114 88092
rect 108941 88090 109007 88093
rect 106108 88088 109007 88090
rect 106108 88032 108946 88088
rect 109002 88032 109007 88088
rect 106108 88030 109007 88032
rect 106108 88028 106114 88030
rect 108941 88027 109007 88030
rect 200062 88028 200068 88092
rect 200132 88090 200138 88092
rect 202505 88090 202571 88093
rect 200132 88088 202571 88090
rect 200132 88032 202510 88088
rect 202566 88032 202571 88088
rect 200132 88030 202571 88032
rect 200132 88028 200138 88030
rect 202505 88027 202571 88030
rect 67909 87818 67975 87821
rect 67909 87816 70380 87818
rect 67909 87760 67914 87816
rect 67970 87760 70380 87816
rect 67909 87758 70380 87760
rect 67909 87755 67975 87758
rect 105670 87756 105676 87820
rect 105740 87756 105746 87820
rect 167085 87818 167151 87821
rect 167085 87816 170292 87818
rect 167085 87760 167090 87816
rect 167146 87760 170292 87816
rect 167085 87758 170292 87760
rect 167085 87755 167151 87758
rect 199694 87756 199700 87820
rect 199764 87756 199770 87820
rect 109769 87546 109835 87549
rect 167678 87546 167684 87548
rect 109769 87544 167684 87546
rect 109769 87488 109774 87544
rect 109830 87488 167684 87544
rect 109769 87486 167684 87488
rect 109769 87483 109835 87486
rect 167678 87484 167684 87486
rect 167748 87546 167754 87548
rect 167748 87486 170322 87546
rect 167748 87484 167754 87486
rect 106038 87348 106044 87412
rect 106108 87410 106114 87412
rect 108481 87410 108547 87413
rect 106108 87408 108547 87410
rect 106108 87352 108486 87408
rect 108542 87352 108547 87408
rect 106108 87350 108547 87352
rect 106108 87348 106114 87350
rect 108481 87347 108547 87350
rect 105670 87076 105676 87140
rect 105740 87076 105746 87140
rect 170262 87108 170322 87486
rect 68093 87002 68159 87005
rect 69289 87002 69355 87005
rect 68093 87000 70380 87002
rect 68093 86944 68098 87000
rect 68154 86944 69294 87000
rect 69350 86944 70380 87000
rect 68093 86942 70380 86944
rect 68093 86939 68159 86942
rect 69289 86939 69355 86942
rect 106038 86668 106044 86732
rect 106108 86730 106114 86732
rect 108941 86730 109007 86733
rect 106108 86728 109007 86730
rect 106108 86672 108946 86728
rect 109002 86672 109007 86728
rect 106108 86670 109007 86672
rect 106108 86668 106114 86670
rect 108941 86667 109007 86670
rect 200062 86668 200068 86732
rect 200132 86730 200138 86732
rect 202505 86730 202571 86733
rect 200132 86728 202571 86730
rect 200132 86672 202510 86728
rect 202566 86672 202571 86728
rect 200132 86670 202571 86672
rect 200132 86668 200138 86670
rect 202505 86667 202571 86670
rect 105670 86396 105676 86460
rect 105740 86396 105746 86460
rect 199694 86396 199700 86460
rect 199764 86396 199770 86460
rect 68829 86322 68895 86325
rect 68829 86320 70380 86322
rect 68829 86264 68834 86320
rect 68890 86264 70380 86320
rect 68829 86262 70380 86264
rect 68829 86259 68895 86262
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 106038 85988 106044 86052
rect 106108 86050 106114 86052
rect 108573 86050 108639 86053
rect 200113 86052 200179 86053
rect 106108 86048 108639 86050
rect 106108 85992 108578 86048
rect 108634 85992 108639 86048
rect 106108 85990 108639 85992
rect 106108 85988 106114 85990
rect 108573 85987 108639 85990
rect 200062 85988 200068 86052
rect 200132 86050 200179 86052
rect 200132 86048 200224 86050
rect 200174 85992 200224 86048
rect 583520 86036 584960 86126
rect 200132 85990 200224 85992
rect 200132 85988 200179 85990
rect 200113 85987 200179 85988
rect 67909 85778 67975 85781
rect 67909 85776 70380 85778
rect 67909 85720 67914 85776
rect 67970 85720 70380 85776
rect 67909 85718 70380 85720
rect 67909 85715 67975 85718
rect 105670 85716 105676 85780
rect 105740 85716 105746 85780
rect 166993 85642 167059 85645
rect 200113 85644 200179 85645
rect 166993 85640 170292 85642
rect 166993 85584 166998 85640
rect 167054 85584 170292 85640
rect 166993 85582 170292 85584
rect 166993 85579 167059 85582
rect 199694 85580 199700 85644
rect 199764 85580 199770 85644
rect 200062 85580 200068 85644
rect 200132 85642 200179 85644
rect 200132 85640 200224 85642
rect 200174 85584 200224 85640
rect 200132 85582 200224 85584
rect 200132 85580 200179 85582
rect 200113 85579 200179 85580
rect 167862 85036 167868 85100
rect 167932 85098 167938 85100
rect 167932 85038 170292 85098
rect 167932 85036 167938 85038
rect 69054 84900 69060 84964
rect 69124 84962 69130 84964
rect 69124 84902 70380 84962
rect 69124 84900 69130 84902
rect 199694 84900 199700 84964
rect 199764 84900 199770 84964
rect -960 84690 480 84780
rect 200062 84764 200068 84828
rect 200132 84826 200138 84828
rect 202689 84826 202755 84829
rect 200132 84824 202755 84826
rect 200132 84768 202694 84824
rect 202750 84768 202755 84824
rect 200132 84766 202755 84768
rect 200132 84764 200138 84766
rect 202689 84763 202755 84766
rect 3417 84690 3483 84693
rect -960 84688 3483 84690
rect -960 84632 3422 84688
rect 3478 84632 3483 84688
rect -960 84630 3483 84632
rect -960 84540 480 84630
rect 3417 84627 3483 84630
rect 106038 84628 106044 84692
rect 106108 84690 106114 84692
rect 108205 84690 108271 84693
rect 106108 84688 108271 84690
rect 106108 84632 108210 84688
rect 108266 84632 108271 84688
rect 106108 84630 108271 84632
rect 106108 84628 106114 84630
rect 108205 84627 108271 84630
rect 67633 84418 67699 84421
rect 67633 84416 70380 84418
rect 67633 84360 67638 84416
rect 67694 84360 70380 84416
rect 67633 84358 70380 84360
rect 67633 84355 67699 84358
rect 105670 84356 105676 84420
rect 105740 84356 105746 84420
rect 167085 84418 167151 84421
rect 167085 84416 170292 84418
rect 167085 84360 167090 84416
rect 167146 84360 170292 84416
rect 167085 84358 170292 84360
rect 167085 84355 167151 84358
rect 199694 84220 199700 84284
rect 199764 84220 199770 84284
rect 200062 84220 200068 84284
rect 200132 84282 200138 84284
rect 202689 84282 202755 84285
rect 200132 84280 202755 84282
rect 200132 84224 202694 84280
rect 202750 84224 202755 84280
rect 200132 84222 202755 84224
rect 200132 84220 200138 84222
rect 202689 84219 202755 84222
rect 106038 83948 106044 84012
rect 106108 84010 106114 84012
rect 108941 84010 109007 84013
rect 106108 84008 109007 84010
rect 106108 83952 108946 84008
rect 109002 83952 109007 84008
rect 106108 83950 109007 83952
rect 106108 83948 106114 83950
rect 108941 83947 109007 83950
rect 105670 83676 105676 83740
rect 105740 83676 105746 83740
rect 66805 83602 66871 83605
rect 68686 83602 68692 83604
rect 66805 83600 68692 83602
rect 66805 83544 66810 83600
rect 66866 83544 68692 83600
rect 66805 83542 68692 83544
rect 66805 83539 66871 83542
rect 68686 83540 68692 83542
rect 68756 83602 68762 83604
rect 68756 83542 70380 83602
rect 68756 83540 68762 83542
rect 106038 83268 106044 83332
rect 106108 83330 106114 83332
rect 109217 83330 109283 83333
rect 170262 83330 170322 83572
rect 199326 83540 199332 83604
rect 199396 83540 199402 83604
rect 106108 83328 109283 83330
rect 106108 83272 109222 83328
rect 109278 83272 109283 83328
rect 106108 83270 109283 83272
rect 106108 83268 106114 83270
rect 109217 83267 109283 83270
rect 113130 83270 170322 83330
rect 106774 83132 106780 83196
rect 106844 83194 106850 83196
rect 113130 83194 113190 83270
rect 200062 83268 200068 83332
rect 200132 83330 200138 83332
rect 203149 83330 203215 83333
rect 200132 83328 203215 83330
rect 200132 83272 203154 83328
rect 203210 83272 203215 83328
rect 200132 83270 203215 83272
rect 200132 83268 200138 83270
rect 203149 83267 203215 83270
rect 106844 83134 113190 83194
rect 106844 83132 106850 83134
rect 105670 82996 105676 83060
rect 105740 82996 105746 83060
rect 166993 83058 167059 83061
rect 166993 83056 170292 83058
rect 166993 83000 166998 83056
rect 167054 83000 170292 83056
rect 166993 82998 170292 83000
rect 166993 82995 167059 82998
rect 199694 82996 199700 83060
rect 199764 82996 199770 83060
rect 200062 82860 200068 82924
rect 200132 82922 200138 82924
rect 201493 82922 201559 82925
rect 200132 82920 201559 82922
rect 200132 82864 201498 82920
rect 201554 82864 201559 82920
rect 200132 82862 201559 82864
rect 200132 82860 200138 82862
rect 201493 82859 201559 82862
rect 106038 82588 106044 82652
rect 106108 82650 106114 82652
rect 108941 82650 109007 82653
rect 106108 82648 109007 82650
rect 106108 82592 108946 82648
rect 109002 82592 109007 82648
rect 106108 82590 109007 82592
rect 106108 82588 106114 82590
rect 108941 82587 109007 82590
rect 105670 82316 105676 82380
rect 105740 82316 105746 82380
rect 69289 82242 69355 82245
rect 69289 82240 70380 82242
rect 69289 82184 69294 82240
rect 69350 82184 70380 82240
rect 69289 82182 70380 82184
rect 69289 82179 69355 82182
rect 106038 81908 106044 81972
rect 106108 81970 106114 81972
rect 108849 81970 108915 81973
rect 170262 81970 170322 82212
rect 199694 82180 199700 82244
rect 199764 82180 199770 82244
rect 106108 81968 108915 81970
rect 106108 81912 108854 81968
rect 108910 81912 108915 81968
rect 106108 81910 108915 81912
rect 106108 81908 106114 81910
rect 108849 81907 108915 81910
rect 113130 81910 170322 81970
rect 106222 81772 106228 81836
rect 106292 81834 106298 81836
rect 113130 81834 113190 81910
rect 200062 81908 200068 81972
rect 200132 81970 200138 81972
rect 202229 81970 202295 81973
rect 200132 81968 202295 81970
rect 200132 81912 202234 81968
rect 202290 81912 202295 81968
rect 200132 81910 202295 81912
rect 200132 81908 200138 81910
rect 202229 81907 202295 81910
rect 106292 81774 113190 81834
rect 106292 81772 106298 81774
rect 105670 81636 105676 81700
rect 105740 81636 105746 81700
rect 68461 81562 68527 81565
rect 166993 81562 167059 81565
rect 68461 81560 70380 81562
rect 68461 81504 68466 81560
rect 68522 81504 70380 81560
rect 68461 81502 70380 81504
rect 166993 81560 170292 81562
rect 166993 81504 166998 81560
rect 167054 81504 170292 81560
rect 166993 81502 170292 81504
rect 68461 81499 68527 81502
rect 166993 81499 167059 81502
rect 106038 81228 106044 81292
rect 106108 81290 106114 81292
rect 108849 81290 108915 81293
rect 106108 81288 108915 81290
rect 106108 81232 108854 81288
rect 108910 81232 108915 81288
rect 106108 81230 108915 81232
rect 106108 81228 106114 81230
rect 108849 81227 108915 81230
rect 105670 80956 105676 81020
rect 105740 80956 105746 81020
rect 67817 80882 67883 80885
rect 68185 80882 68251 80885
rect 67817 80880 70380 80882
rect 67817 80824 67822 80880
rect 67878 80824 68190 80880
rect 68246 80824 70380 80880
rect 67817 80822 70380 80824
rect 67817 80819 67883 80822
rect 68185 80819 68251 80822
rect 199694 80820 199700 80884
rect 199764 80820 199770 80884
rect 106038 80548 106044 80612
rect 106108 80610 106114 80612
rect 108941 80610 109007 80613
rect 106108 80608 109007 80610
rect 106108 80552 108946 80608
rect 109002 80552 109007 80608
rect 106108 80550 109007 80552
rect 106108 80548 106114 80550
rect 108941 80547 109007 80550
rect 200062 80548 200068 80612
rect 200132 80610 200138 80612
rect 202045 80610 202111 80613
rect 200132 80608 202111 80610
rect 200132 80552 202050 80608
rect 202106 80552 202111 80608
rect 200132 80550 202111 80552
rect 200132 80548 200138 80550
rect 202045 80547 202111 80550
rect 105670 80276 105676 80340
rect 105740 80276 105746 80340
rect 166993 80338 167059 80341
rect 166993 80336 170292 80338
rect 166993 80280 166998 80336
rect 167054 80280 170292 80336
rect 166993 80278 170292 80280
rect 166993 80275 167059 80278
rect 69749 80202 69815 80205
rect 69749 80200 70380 80202
rect 69749 80144 69754 80200
rect 69810 80144 70380 80200
rect 69749 80142 70380 80144
rect 69749 80139 69815 80142
rect 199694 80140 199700 80204
rect 199764 80140 199770 80204
rect 202505 80202 202571 80205
rect 200070 80200 202571 80202
rect 200070 80144 202510 80200
rect 202566 80144 202571 80200
rect 200070 80142 202571 80144
rect 200070 80068 200130 80142
rect 202505 80139 202571 80142
rect 200062 80004 200068 80068
rect 200132 80004 200138 80068
rect 106038 79868 106044 79932
rect 106108 79930 106114 79932
rect 107745 79930 107811 79933
rect 106108 79928 107811 79930
rect 106108 79872 107750 79928
rect 107806 79872 107811 79928
rect 106108 79870 107811 79872
rect 106108 79868 106114 79870
rect 107745 79867 107811 79870
rect 105670 79596 105676 79660
rect 105740 79596 105746 79660
rect 69381 79522 69447 79525
rect 167637 79522 167703 79525
rect 168281 79522 168347 79525
rect 69381 79520 70380 79522
rect 69381 79464 69386 79520
rect 69442 79464 70380 79520
rect 69381 79462 70380 79464
rect 167637 79520 170292 79522
rect 167637 79464 167642 79520
rect 167698 79464 168286 79520
rect 168342 79464 170292 79520
rect 167637 79462 170292 79464
rect 69381 79459 69447 79462
rect 167637 79459 167703 79462
rect 168281 79459 168347 79462
rect 199694 79460 199700 79524
rect 199764 79460 199770 79524
rect 106038 79188 106044 79252
rect 106108 79250 106114 79252
rect 108665 79250 108731 79253
rect 106108 79248 108731 79250
rect 106108 79192 108670 79248
rect 108726 79192 108731 79248
rect 106108 79190 108731 79192
rect 106108 79188 106114 79190
rect 108665 79187 108731 79190
rect 200062 79188 200068 79252
rect 200132 79250 200138 79252
rect 202781 79250 202847 79253
rect 200132 79248 202847 79250
rect 200132 79192 202786 79248
rect 202842 79192 202847 79248
rect 200132 79190 202847 79192
rect 200132 79188 200138 79190
rect 202781 79187 202847 79190
rect 105670 78916 105676 78980
rect 105740 78916 105746 78980
rect 67633 78842 67699 78845
rect 68001 78842 68067 78845
rect 166993 78842 167059 78845
rect 67633 78840 70380 78842
rect 67633 78784 67638 78840
rect 67694 78784 68006 78840
rect 68062 78784 70380 78840
rect 67633 78782 70380 78784
rect 166993 78840 170292 78842
rect 166993 78784 166998 78840
rect 167054 78784 170292 78840
rect 166993 78782 170292 78784
rect 67633 78779 67699 78782
rect 68001 78779 68067 78782
rect 166993 78779 167059 78782
rect 199694 78780 199700 78844
rect 199764 78780 199770 78844
rect 200062 78644 200068 78708
rect 200132 78706 200138 78708
rect 202781 78706 202847 78709
rect 200132 78704 202847 78706
rect 200132 78648 202786 78704
rect 202842 78648 202847 78704
rect 200132 78646 202847 78648
rect 200132 78644 200138 78646
rect 202781 78643 202847 78646
rect 67633 78298 67699 78301
rect 67633 78296 70380 78298
rect 67633 78240 67638 78296
rect 67694 78240 70380 78296
rect 67633 78238 70380 78240
rect 67633 78235 67699 78238
rect 167729 78162 167795 78165
rect 167729 78160 170292 78162
rect 167729 78104 167734 78160
rect 167790 78104 170292 78160
rect 167729 78102 170292 78104
rect 167729 78099 167795 78102
rect 199326 78100 199332 78164
rect 199396 78100 199402 78164
rect 106038 77828 106044 77892
rect 106108 77890 106114 77892
rect 107745 77890 107811 77893
rect 106108 77888 107811 77890
rect 106108 77832 107750 77888
rect 107806 77832 107811 77888
rect 106108 77830 107811 77832
rect 106108 77828 106114 77830
rect 107745 77827 107811 77830
rect 67633 77618 67699 77621
rect 67633 77616 70380 77618
rect 67633 77560 67638 77616
rect 67694 77560 70380 77616
rect 67633 77558 70380 77560
rect 67633 77555 67699 77558
rect 105670 77556 105676 77620
rect 105740 77556 105746 77620
rect 168281 77482 168347 77485
rect 168281 77480 170292 77482
rect 168281 77424 168286 77480
rect 168342 77424 170292 77480
rect 168281 77422 170292 77424
rect 168281 77419 168347 77422
rect 199694 77420 199700 77484
rect 199764 77420 199770 77484
rect 200062 77284 200068 77348
rect 200132 77346 200138 77348
rect 200665 77346 200731 77349
rect 200132 77344 200731 77346
rect 200132 77288 200670 77344
rect 200726 77288 200731 77344
rect 200132 77286 200731 77288
rect 200132 77284 200138 77286
rect 200665 77283 200731 77286
rect 106181 77210 106247 77213
rect 107745 77210 107811 77213
rect 106181 77208 107811 77210
rect 106181 77152 106186 77208
rect 106242 77152 107750 77208
rect 107806 77152 107811 77208
rect 106181 77150 107811 77152
rect 106181 77147 106247 77150
rect 107745 77147 107811 77150
rect 168189 76938 168255 76941
rect 168189 76936 170292 76938
rect 168189 76880 168194 76936
rect 168250 76880 170292 76936
rect 168189 76878 170292 76880
rect 168189 76875 168255 76878
rect 69473 76802 69539 76805
rect 69473 76800 70380 76802
rect 69473 76744 69478 76800
rect 69534 76744 70380 76800
rect 69473 76742 70380 76744
rect 69473 76739 69539 76742
rect 105670 76740 105676 76804
rect 105740 76740 105746 76804
rect 199694 76740 199700 76804
rect 199764 76740 199770 76804
rect 106038 76468 106044 76532
rect 106108 76530 106114 76532
rect 106181 76530 106247 76533
rect 106108 76528 106247 76530
rect 106108 76472 106186 76528
rect 106242 76472 106247 76528
rect 106108 76470 106247 76472
rect 106108 76468 106114 76470
rect 106181 76467 106247 76470
rect 106406 76468 106412 76532
rect 106476 76530 106482 76532
rect 106476 76470 170322 76530
rect 106476 76468 106482 76470
rect 170262 76228 170322 76470
rect 200062 76468 200068 76532
rect 200132 76530 200138 76532
rect 201309 76530 201375 76533
rect 200132 76528 201375 76530
rect 200132 76472 201314 76528
rect 201370 76472 201375 76528
rect 200132 76470 201375 76472
rect 200132 76468 200138 76470
rect 201309 76467 201375 76470
rect 105670 76060 105676 76124
rect 105740 76060 105746 76124
rect 106038 75924 106044 75988
rect 106108 75986 106114 75988
rect 107745 75986 107811 75989
rect 106108 75984 107811 75986
rect 106108 75928 107750 75984
rect 107806 75928 107811 75984
rect 106108 75926 107811 75928
rect 106108 75924 106114 75926
rect 107745 75923 107811 75926
rect 67725 75850 67791 75853
rect 68921 75850 68987 75853
rect 107837 75850 107903 75853
rect 67725 75848 68987 75850
rect 67725 75792 67730 75848
rect 67786 75792 68926 75848
rect 68982 75792 68987 75848
rect 67725 75790 68987 75792
rect 67725 75787 67791 75790
rect 68921 75787 68987 75790
rect 106046 75848 107903 75850
rect 106046 75792 107842 75848
rect 107898 75792 107903 75848
rect 106046 75790 107903 75792
rect 106046 75716 106106 75790
rect 107837 75787 107903 75790
rect 67398 75652 67404 75716
rect 67468 75714 67474 75716
rect 68870 75714 68876 75716
rect 67468 75654 68876 75714
rect 67468 75652 67474 75654
rect 68870 75652 68876 75654
rect 68940 75652 68946 75716
rect 106038 75652 106044 75716
rect 106108 75652 106114 75716
rect 68878 75578 68938 75652
rect 68878 75518 70380 75578
rect 105670 75516 105676 75580
rect 105740 75516 105746 75580
rect 199694 75380 199700 75444
rect 199764 75380 199770 75444
rect 106038 75108 106044 75172
rect 106108 75170 106114 75172
rect 107745 75170 107811 75173
rect 106108 75168 107811 75170
rect 106108 75112 107750 75168
rect 107806 75112 107811 75168
rect 106108 75110 107811 75112
rect 106108 75108 106114 75110
rect 107745 75107 107811 75110
rect 200062 75108 200068 75172
rect 200132 75170 200138 75172
rect 200481 75170 200547 75173
rect 200132 75168 200547 75170
rect 200132 75112 200486 75168
rect 200542 75112 200547 75168
rect 200132 75110 200547 75112
rect 200132 75108 200138 75110
rect 200481 75107 200547 75110
rect 106181 75036 106247 75037
rect 106181 75034 106228 75036
rect 106136 75032 106228 75034
rect 106136 74976 106186 75032
rect 106136 74974 106228 74976
rect 106181 74972 106228 74974
rect 106292 74972 106298 75036
rect 106181 74971 106247 74972
rect 68921 74898 68987 74901
rect 68921 74896 70380 74898
rect 68921 74840 68926 74896
rect 68982 74840 70380 74896
rect 68921 74838 70380 74840
rect 68921 74835 68987 74838
rect 105670 74836 105676 74900
rect 105740 74836 105746 74900
rect 167085 74762 167151 74765
rect 167085 74760 170292 74762
rect 167085 74704 167090 74760
rect 167146 74704 170292 74760
rect 167085 74702 170292 74704
rect 167085 74699 167151 74702
rect 199326 74700 199332 74764
rect 199396 74700 199402 74764
rect 200062 74700 200068 74764
rect 200132 74762 200138 74764
rect 200941 74762 201007 74765
rect 200132 74760 201007 74762
rect 200132 74704 200946 74760
rect 201002 74704 201007 74760
rect 200132 74702 201007 74704
rect 200132 74700 200138 74702
rect 200941 74699 201007 74702
rect 107745 74490 107811 74493
rect 106046 74488 107811 74490
rect 106046 74432 107750 74488
rect 107806 74432 107811 74488
rect 106046 74430 107811 74432
rect 68502 74020 68508 74084
rect 68572 74082 68578 74084
rect 68829 74082 68895 74085
rect 106046 74084 106106 74430
rect 107745 74427 107811 74430
rect 68572 74080 70380 74082
rect 68572 74024 68834 74080
rect 68890 74024 70380 74080
rect 68572 74022 70380 74024
rect 68572 74020 68578 74022
rect 68829 74019 68895 74022
rect 105670 74020 105676 74084
rect 105740 74020 105746 74084
rect 106038 74020 106044 74084
rect 106108 74020 106114 74084
rect 167085 74082 167151 74085
rect 167085 74080 170292 74082
rect 167085 74024 167090 74080
rect 167146 74024 170292 74080
rect 167085 74022 170292 74024
rect 167085 74019 167151 74022
rect 199694 74020 199700 74084
rect 199764 74020 199770 74084
rect 153101 73946 153167 73949
rect 168966 73946 168972 73948
rect 153101 73944 168972 73946
rect 153101 73888 153106 73944
rect 153162 73888 168972 73944
rect 153101 73886 168972 73888
rect 153101 73883 153167 73886
rect 168966 73884 168972 73886
rect 169036 73884 169042 73948
rect 113081 73810 113147 73813
rect 170254 73810 170260 73812
rect 106046 73808 170260 73810
rect 106046 73752 113086 73808
rect 113142 73752 170260 73808
rect 106046 73750 170260 73752
rect 106046 73676 106106 73750
rect 113081 73747 113147 73750
rect 170254 73748 170260 73750
rect 170324 73748 170330 73812
rect 200062 73748 200068 73812
rect 200132 73810 200138 73812
rect 200849 73810 200915 73813
rect 201953 73810 202019 73813
rect 200132 73808 202019 73810
rect 200132 73752 200854 73808
rect 200910 73752 201958 73808
rect 202014 73752 202019 73808
rect 200132 73750 202019 73752
rect 200132 73748 200138 73750
rect 200849 73747 200915 73750
rect 201953 73747 202019 73750
rect 106038 73612 106044 73676
rect 106108 73612 106114 73676
rect 69238 73340 69244 73404
rect 69308 73402 69314 73404
rect 69308 73372 70564 73402
rect 69308 73342 70594 73372
rect 69308 73340 69314 73342
rect 68318 73204 68324 73268
rect 68388 73266 68394 73268
rect 69565 73266 69631 73269
rect 70534 73268 70594 73342
rect 105670 73340 105676 73404
rect 105740 73340 105746 73404
rect 167177 73402 167243 73405
rect 167177 73400 170292 73402
rect 167177 73344 167182 73400
rect 167238 73344 170292 73400
rect 167177 73342 170292 73344
rect 167177 73339 167243 73342
rect 199694 73340 199700 73404
rect 199764 73340 199770 73404
rect 68388 73264 69631 73266
rect 68388 73208 69570 73264
rect 69626 73208 69631 73264
rect 68388 73206 69631 73208
rect 68388 73204 68394 73206
rect 69565 73203 69631 73206
rect 70526 73204 70532 73268
rect 70596 73204 70602 73268
rect 200062 73204 200068 73268
rect 200132 73266 200138 73268
rect 200573 73266 200639 73269
rect 200132 73264 200639 73266
rect 200132 73208 200578 73264
rect 200634 73208 200639 73264
rect 200132 73206 200639 73208
rect 200132 73204 200138 73206
rect 200573 73203 200639 73206
rect 107837 73130 107903 73133
rect 106046 73128 107903 73130
rect 106046 73072 107842 73128
rect 107898 73072 107903 73128
rect 106046 73070 107903 73072
rect 106046 72860 106106 73070
rect 107837 73067 107903 73070
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 106038 72796 106044 72860
rect 106108 72796 106114 72860
rect 583520 72844 584960 72934
rect 69565 72722 69631 72725
rect 69565 72720 70380 72722
rect 69565 72664 69570 72720
rect 69626 72664 70380 72720
rect 69565 72662 70380 72664
rect 69565 72659 69631 72662
rect 105670 72660 105676 72724
rect 105740 72660 105746 72724
rect 167862 72660 167868 72724
rect 167932 72722 167938 72724
rect 167932 72662 170292 72722
rect 167932 72660 167938 72662
rect 199694 72660 199700 72724
rect 199764 72660 199770 72724
rect 107745 72450 107811 72453
rect 106046 72448 107811 72450
rect 106046 72392 107750 72448
rect 107806 72392 107811 72448
rect 106046 72390 107811 72392
rect 106046 72316 106106 72390
rect 107745 72387 107811 72390
rect 200062 72388 200068 72452
rect 200132 72450 200138 72452
rect 200757 72450 200823 72453
rect 200132 72448 200823 72450
rect 200132 72392 200762 72448
rect 200818 72392 200823 72448
rect 200132 72390 200823 72392
rect 200132 72388 200138 72390
rect 200757 72387 200823 72390
rect 106038 72252 106044 72316
rect 106108 72252 106114 72316
rect 105670 72116 105676 72180
rect 105740 72116 105746 72180
rect 68277 72042 68343 72045
rect 167085 72042 167151 72045
rect 68277 72040 70380 72042
rect 68277 71984 68282 72040
rect 68338 71984 70380 72040
rect 68277 71982 70380 71984
rect 167085 72040 170292 72042
rect 167085 71984 167090 72040
rect 167146 71984 170292 72040
rect 167085 71982 170292 71984
rect 68277 71979 68343 71982
rect 167085 71979 167151 71982
rect 199694 71980 199700 72044
rect 199764 71980 199770 72044
rect 200062 71844 200068 71908
rect 200132 71906 200138 71908
rect 200205 71906 200271 71909
rect 200132 71904 200271 71906
rect 200132 71848 200210 71904
rect 200266 71848 200271 71904
rect 200132 71846 200271 71848
rect 200132 71844 200138 71846
rect 200205 71843 200271 71846
rect -960 71634 480 71724
rect 2865 71634 2931 71637
rect -960 71632 2931 71634
rect -960 71576 2870 71632
rect 2926 71576 2931 71632
rect -960 71574 2931 71576
rect -960 71484 480 71574
rect 2865 71571 2931 71574
rect 68645 71362 68711 71365
rect 69841 71362 69907 71365
rect 168005 71362 168071 71365
rect 68645 71360 70380 71362
rect 68645 71304 68650 71360
rect 68706 71304 69846 71360
rect 69902 71304 70380 71360
rect 68645 71302 70380 71304
rect 168005 71360 170292 71362
rect 168005 71304 168010 71360
rect 168066 71304 170292 71360
rect 168005 71302 170292 71304
rect 68645 71299 68711 71302
rect 69841 71299 69907 71302
rect 168005 71299 168071 71302
rect 199702 71226 199762 71332
rect 201953 71226 202019 71229
rect 199702 71224 202019 71226
rect 199702 71168 201958 71224
rect 202014 71168 202019 71224
rect 199702 71166 202019 71168
rect 106038 71028 106044 71092
rect 106108 71090 106114 71092
rect 113081 71090 113147 71093
rect 116577 71090 116643 71093
rect 106108 71088 116643 71090
rect 106108 71032 113086 71088
rect 113142 71032 116582 71088
rect 116638 71032 116643 71088
rect 106108 71030 116643 71032
rect 106108 71028 106114 71030
rect 113081 71027 113147 71030
rect 116577 71027 116643 71030
rect 69657 70682 69723 70685
rect 69657 70680 70380 70682
rect 69657 70624 69662 70680
rect 69718 70624 70380 70680
rect 69657 70622 70380 70624
rect 69657 70619 69723 70622
rect 105670 70620 105676 70684
rect 105740 70620 105746 70684
rect 168097 70682 168163 70685
rect 198733 70682 198799 70685
rect 199702 70682 199762 71166
rect 201953 71163 202019 71166
rect 168097 70680 170292 70682
rect 168097 70624 168102 70680
rect 168158 70624 170292 70680
rect 168097 70622 170292 70624
rect 198733 70680 199762 70682
rect 198733 70624 198738 70680
rect 198794 70624 199762 70680
rect 198733 70622 199762 70624
rect 168097 70619 168163 70622
rect 198733 70619 198799 70622
rect 202045 70546 202111 70549
rect 195930 70544 202111 70546
rect 195930 70488 202050 70544
rect 202106 70488 202111 70544
rect 195930 70486 202111 70488
rect 106181 70410 106247 70413
rect 106046 70408 106247 70410
rect 106046 70352 106186 70408
rect 106242 70352 106247 70408
rect 106046 70350 106247 70352
rect 106046 70276 106106 70350
rect 106181 70347 106247 70350
rect 167453 70410 167519 70413
rect 170029 70410 170095 70413
rect 195930 70410 195990 70486
rect 202045 70483 202111 70486
rect 167453 70408 170095 70410
rect 167453 70352 167458 70408
rect 167514 70352 170034 70408
rect 170090 70352 170095 70408
rect 167453 70350 170095 70352
rect 167453 70347 167519 70350
rect 170029 70347 170095 70350
rect 180750 70350 195990 70410
rect 106038 70212 106044 70276
rect 106108 70212 106114 70276
rect 105670 70076 105676 70140
rect 105740 70076 105746 70140
rect 70301 70002 70367 70005
rect 70526 70002 70532 70004
rect 70301 70000 70532 70002
rect 70301 69944 70306 70000
rect 70362 69944 70532 70000
rect 70301 69942 70532 69944
rect 70301 69939 70367 69942
rect 70526 69940 70532 69942
rect 70596 69940 70602 70004
rect 69054 69804 69060 69868
rect 69124 69866 69130 69868
rect 167678 69866 167684 69868
rect 69124 69806 167684 69866
rect 69124 69804 69130 69806
rect 167678 69804 167684 69806
rect 167748 69804 167754 69868
rect 168966 69804 168972 69868
rect 169036 69866 169042 69868
rect 180750 69866 180810 70350
rect 169036 69806 180810 69866
rect 199334 69869 199394 69972
rect 199334 69864 199443 69869
rect 199334 69808 199382 69864
rect 199438 69808 199443 69864
rect 199334 69806 199443 69808
rect 169036 69804 169042 69806
rect 199377 69803 199443 69806
rect 69197 69730 69263 69733
rect 167310 69730 167316 69732
rect 69197 69728 167316 69730
rect 69197 69672 69202 69728
rect 69258 69672 167316 69728
rect 69197 69670 167316 69672
rect 69197 69667 69263 69670
rect 167310 69668 167316 69670
rect 167380 69668 167386 69732
rect 170254 69668 170260 69732
rect 170324 69730 170330 69732
rect 202505 69730 202571 69733
rect 170324 69728 202571 69730
rect 170324 69672 202510 69728
rect 202566 69672 202571 69728
rect 170324 69670 202571 69672
rect 170324 69668 170330 69670
rect 202505 69667 202571 69670
rect 68686 69532 68692 69596
rect 68756 69594 68762 69596
rect 106774 69594 106780 69596
rect 68756 69534 106780 69594
rect 68756 69532 68762 69534
rect 106774 69532 106780 69534
rect 106844 69532 106850 69596
rect 166809 69594 166875 69597
rect 201718 69594 201724 69596
rect 166809 69592 201724 69594
rect 166809 69536 166814 69592
rect 166870 69536 201724 69592
rect 166809 69534 201724 69536
rect 166809 69531 166875 69534
rect 201718 69532 201724 69534
rect 201788 69532 201794 69596
rect 68870 69396 68876 69460
rect 68940 69458 68946 69460
rect 106038 69458 106044 69460
rect 68940 69398 106044 69458
rect 68940 69396 68946 69398
rect 106038 69396 106044 69398
rect 106108 69396 106114 69460
rect 113541 69458 113607 69461
rect 199326 69458 199332 69460
rect 113541 69456 199332 69458
rect 113541 69400 113546 69456
rect 113602 69400 199332 69456
rect 113541 69398 199332 69400
rect 113541 69395 113607 69398
rect 199326 69396 199332 69398
rect 199396 69396 199402 69460
rect 105486 69260 105492 69324
rect 105556 69322 105562 69324
rect 113817 69322 113883 69325
rect 199142 69322 199148 69324
rect 105556 69320 199148 69322
rect 105556 69264 113822 69320
rect 113878 69264 199148 69320
rect 105556 69262 199148 69264
rect 105556 69260 105562 69262
rect 113817 69259 113883 69262
rect 199142 69260 199148 69262
rect 199212 69260 199218 69324
rect 89345 68914 89411 68917
rect 115933 68914 115999 68917
rect 117221 68914 117287 68917
rect 89345 68912 117287 68914
rect 89345 68856 89350 68912
rect 89406 68856 115938 68912
rect 115994 68856 117226 68912
rect 117282 68856 117287 68912
rect 89345 68854 117287 68856
rect 89345 68851 89411 68854
rect 115933 68851 115999 68854
rect 117221 68851 117287 68854
rect 163405 68914 163471 68917
rect 164049 68914 164115 68917
rect 171317 68914 171383 68917
rect 171869 68914 171935 68917
rect 163405 68912 171935 68914
rect 163405 68856 163410 68912
rect 163466 68856 164054 68912
rect 164110 68856 171322 68912
rect 171378 68856 171874 68912
rect 171930 68856 171935 68912
rect 163405 68854 171935 68856
rect 163405 68851 163471 68854
rect 164049 68851 164115 68854
rect 171317 68851 171383 68854
rect 171869 68851 171935 68854
rect 189073 68914 189139 68917
rect 190361 68914 190427 68917
rect 200062 68914 200068 68916
rect 189073 68912 200068 68914
rect 189073 68856 189078 68912
rect 189134 68856 190366 68912
rect 190422 68856 200068 68912
rect 189073 68854 200068 68856
rect 189073 68851 189139 68854
rect 190361 68851 190427 68854
rect 200062 68852 200068 68854
rect 200132 68852 200138 68916
rect 77753 68778 77819 68781
rect 163865 68778 163931 68781
rect 177297 68778 177363 68781
rect 177757 68778 177823 68781
rect 77753 68776 177823 68778
rect 77753 68720 77758 68776
rect 77814 68720 163870 68776
rect 163926 68720 177302 68776
rect 177358 68720 177762 68776
rect 177818 68720 177823 68776
rect 77753 68718 177823 68720
rect 77753 68715 77819 68718
rect 163865 68715 163931 68718
rect 177297 68715 177363 68718
rect 177757 68715 177823 68718
rect 95141 68642 95207 68645
rect 113357 68642 113423 68645
rect 192569 68642 192635 68645
rect 95141 68640 192635 68642
rect 95141 68584 95146 68640
rect 95202 68584 113362 68640
rect 113418 68584 192574 68640
rect 192630 68584 192635 68640
rect 95141 68582 192635 68584
rect 95141 68579 95207 68582
rect 113357 68579 113423 68582
rect 192569 68579 192635 68582
rect 84193 68506 84259 68509
rect 114645 68506 114711 68509
rect 115841 68506 115907 68509
rect 84193 68504 115907 68506
rect 84193 68448 84198 68504
rect 84254 68448 114650 68504
rect 114706 68448 115846 68504
rect 115902 68448 115907 68504
rect 84193 68446 115907 68448
rect 84193 68443 84259 68446
rect 114645 68443 114711 68446
rect 115841 68443 115907 68446
rect 117221 68506 117287 68509
rect 189073 68506 189139 68509
rect 117221 68504 189139 68506
rect 117221 68448 117226 68504
rect 117282 68448 189078 68504
rect 189134 68448 189139 68504
rect 117221 68446 189139 68448
rect 117221 68443 117287 68446
rect 189073 68443 189139 68446
rect 79685 68370 79751 68373
rect 116669 68370 116735 68373
rect 179689 68370 179755 68373
rect 180057 68370 180123 68373
rect 79685 68368 180123 68370
rect 79685 68312 79690 68368
rect 79746 68312 116674 68368
rect 116730 68312 179694 68368
rect 179750 68312 180062 68368
rect 180118 68312 180123 68368
rect 79685 68310 180123 68312
rect 79685 68307 79751 68310
rect 116669 68307 116735 68310
rect 179689 68307 179755 68310
rect 180057 68307 180123 68310
rect 74533 68234 74599 68237
rect 111241 68234 111307 68237
rect 174537 68234 174603 68237
rect 74533 68232 174603 68234
rect 74533 68176 74538 68232
rect 74594 68176 111246 68232
rect 111302 68176 174542 68232
rect 174598 68176 174603 68232
rect 74533 68174 174603 68176
rect 74533 68171 74599 68174
rect 111241 68171 111307 68174
rect 174537 68171 174603 68174
rect 115841 68098 115907 68101
rect 166257 68098 166323 68101
rect 115841 68096 166323 68098
rect 115841 68040 115846 68096
rect 115902 68040 166262 68096
rect 166318 68040 166323 68096
rect 115841 68038 166323 68040
rect 115841 68035 115907 68038
rect 166257 68035 166323 68038
rect 70393 67962 70459 67965
rect 163405 67962 163471 67965
rect 70393 67960 163471 67962
rect 70393 67904 70398 67960
rect 70454 67904 163410 67960
rect 163466 67904 163471 67960
rect 70393 67902 163471 67904
rect 70393 67899 70459 67902
rect 163405 67899 163471 67902
rect 165337 67554 165403 67557
rect 165521 67554 165587 67557
rect 188705 67554 188771 67557
rect 165337 67552 188771 67554
rect 165337 67496 165342 67552
rect 165398 67496 165526 67552
rect 165582 67496 188710 67552
rect 188766 67496 188771 67552
rect 165337 67494 188771 67496
rect 165337 67491 165403 67494
rect 165521 67491 165587 67494
rect 188705 67491 188771 67494
rect 100937 67418 101003 67421
rect 141509 67418 141575 67421
rect 200205 67418 200271 67421
rect 100937 67416 200271 67418
rect 100937 67360 100942 67416
rect 100998 67360 141514 67416
rect 141570 67360 200210 67416
rect 200266 67360 200271 67416
rect 100937 67358 200271 67360
rect 100937 67355 101003 67358
rect 141509 67355 141575 67358
rect 200205 67355 200271 67358
rect 68461 67282 68527 67285
rect 105302 67282 105308 67284
rect 68461 67280 105308 67282
rect 68461 67224 68466 67280
rect 68522 67224 105308 67280
rect 68461 67222 105308 67224
rect 68461 67219 68527 67222
rect 105302 67220 105308 67222
rect 105372 67220 105378 67284
rect 166349 67282 166415 67285
rect 201534 67282 201540 67284
rect 166349 67280 201540 67282
rect 166349 67224 166354 67280
rect 166410 67224 201540 67280
rect 166349 67222 201540 67224
rect 166349 67219 166415 67222
rect 201534 67220 201540 67222
rect 201604 67220 201610 67284
rect 88057 67146 88123 67149
rect 165521 67146 165587 67149
rect 88057 67144 165587 67146
rect 88057 67088 88062 67144
rect 88118 67088 165526 67144
rect 165582 67088 165587 67144
rect 88057 67086 165587 67088
rect 88057 67083 88123 67086
rect 165521 67083 165587 67086
rect 103513 66194 103579 66197
rect 200849 66194 200915 66197
rect 103513 66192 200915 66194
rect 103513 66136 103518 66192
rect 103574 66136 200854 66192
rect 200910 66136 200915 66192
rect 103513 66134 200915 66136
rect 103513 66131 103579 66134
rect 200849 66131 200915 66134
rect 106273 66058 106339 66061
rect 107009 66058 107075 66061
rect 173249 66058 173315 66061
rect 106273 66056 173315 66058
rect 106273 66000 106278 66056
rect 106334 66000 107014 66056
rect 107070 66000 173254 66056
rect 173310 66000 173315 66056
rect 106273 65998 173315 66000
rect 106273 65995 106339 65998
rect 107009 65995 107075 65998
rect 173249 65995 173315 65998
rect 78397 65922 78463 65925
rect 113909 65922 113975 65925
rect 178401 65922 178467 65925
rect 78397 65920 178467 65922
rect 78397 65864 78402 65920
rect 78458 65864 113914 65920
rect 113970 65864 178406 65920
rect 178462 65864 178467 65920
rect 78397 65862 178467 65864
rect 78397 65859 78463 65862
rect 113909 65859 113975 65862
rect 178401 65859 178467 65862
rect 68277 65786 68343 65789
rect 107561 65786 107627 65789
rect 68277 65784 107627 65786
rect 68277 65728 68282 65784
rect 68338 65728 107566 65784
rect 107622 65728 107627 65784
rect 68277 65726 107627 65728
rect 68277 65723 68343 65726
rect 107561 65723 107627 65726
rect 69565 64834 69631 64837
rect 167862 64834 167868 64836
rect 69565 64832 167868 64834
rect 69565 64776 69570 64832
rect 69626 64776 167868 64832
rect 69565 64774 167868 64776
rect 69565 64771 69631 64774
rect 167862 64772 167868 64774
rect 167932 64772 167938 64836
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3509 58578 3575 58581
rect -960 58576 3575 58578
rect -960 58520 3514 58576
rect 3570 58520 3575 58576
rect -960 58518 3575 58520
rect -960 58428 480 58518
rect 3509 58515 3575 58518
rect 167862 58516 167868 58580
rect 167932 58578 167938 58580
rect 328453 58578 328519 58581
rect 167932 58576 328519 58578
rect 167932 58520 328458 58576
rect 328514 58520 328519 58576
rect 167932 58518 328519 58520
rect 167932 58516 167938 58518
rect 328453 58515 328519 58518
rect 170070 57156 170076 57220
rect 170140 57218 170146 57220
rect 309133 57218 309199 57221
rect 170140 57216 309199 57218
rect 170140 57160 309138 57216
rect 309194 57160 309199 57216
rect 170140 57158 309199 57160
rect 170140 57156 170146 57158
rect 309133 57155 309199 57158
rect 167494 54436 167500 54500
rect 167564 54498 167570 54500
rect 338113 54498 338179 54501
rect 167564 54496 338179 54498
rect 167564 54440 338118 54496
rect 338174 54440 338179 54496
rect 167564 54438 338179 54440
rect 167564 54436 167570 54438
rect 338113 54435 338179 54438
rect 169334 53076 169340 53140
rect 169404 53138 169410 53140
rect 340965 53138 341031 53141
rect 169404 53136 341031 53138
rect 169404 53080 340970 53136
rect 341026 53080 341031 53136
rect 169404 53078 341031 53080
rect 169404 53076 169410 53078
rect 340965 53075 341031 53078
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 2773 45522 2839 45525
rect -960 45520 2839 45522
rect -960 45464 2778 45520
rect 2834 45464 2839 45520
rect -960 45462 2839 45464
rect -960 45372 480 45462
rect 2773 45459 2839 45462
rect 169702 43420 169708 43484
rect 169772 43482 169778 43484
rect 303613 43482 303679 43485
rect 169772 43480 303679 43482
rect 169772 43424 303618 43480
rect 303674 43424 303679 43480
rect 169772 43422 303679 43424
rect 169772 43420 169778 43422
rect 303613 43419 303679 43422
rect 169886 40564 169892 40628
rect 169956 40626 169962 40628
rect 335353 40626 335419 40629
rect 169956 40624 335419 40626
rect 169956 40568 335358 40624
rect 335414 40568 335419 40624
rect 169956 40566 335419 40568
rect 169956 40564 169962 40566
rect 335353 40563 335419 40566
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2865 32466 2931 32469
rect -960 32464 2931 32466
rect -960 32408 2870 32464
rect 2926 32408 2931 32464
rect -960 32406 2931 32408
rect -960 32316 480 32406
rect 2865 32403 2931 32406
rect 169518 19892 169524 19956
rect 169588 19954 169594 19956
rect 332685 19954 332751 19957
rect 169588 19952 332751 19954
rect 169588 19896 332690 19952
rect 332746 19896 332751 19952
rect 169588 19894 332751 19896
rect 169588 19892 169594 19894
rect 332685 19891 332751 19894
rect 580257 19818 580323 19821
rect 583520 19818 584960 19908
rect 580257 19816 584960 19818
rect 580257 19760 580262 19816
rect 580318 19760 584960 19816
rect 580257 19758 584960 19760
rect 580257 19755 580323 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3509 19410 3575 19413
rect -960 19408 3575 19410
rect -960 19352 3514 19408
rect 3570 19352 3575 19408
rect -960 19350 3575 19352
rect -960 19260 480 19350
rect 3509 19347 3575 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< via3 >>
rect 68324 252860 68388 252924
rect 68692 252724 68756 252788
rect 68508 252588 68572 252652
rect 120028 251908 120092 251972
rect 69060 251772 69124 251836
rect 119844 251500 119908 251564
rect 119476 250140 119540 250204
rect 119660 250004 119724 250068
rect 68876 248296 68940 248300
rect 68876 248240 68890 248296
rect 68890 248240 68940 248296
rect 68876 248236 68940 248240
rect 119844 247964 119908 248028
rect 120028 247556 120092 247620
rect 121868 246196 121932 246260
rect 122236 242992 122300 242996
rect 122236 242936 122286 242992
rect 122286 242936 122300 242992
rect 122236 242932 122300 242936
rect 67220 241572 67284 241636
rect 120212 240212 120276 240276
rect 230428 240212 230492 240276
rect 68324 239532 68388 239596
rect 68508 238852 68572 238916
rect 169524 233820 169588 233884
rect 119844 233004 119908 233068
rect 68692 232656 68756 232660
rect 68692 232600 68742 232656
rect 68742 232600 68756 232656
rect 68692 232596 68756 232600
rect 119476 232460 119540 232524
rect 169708 230556 169772 230620
rect 119660 229196 119724 229260
rect 119292 228516 119356 228580
rect 120028 227836 120092 227900
rect 231900 227700 231964 227764
rect 120580 226340 120644 226404
rect 119292 221172 119356 221236
rect 167500 217636 167564 217700
rect 230428 217908 230492 217972
rect 122052 213012 122116 213076
rect 119292 210700 119356 210764
rect 68692 210156 68756 210220
rect 122420 210156 122484 210220
rect 70716 209476 70780 209540
rect 69244 207436 69308 207500
rect 68508 205532 68572 205596
rect 69796 204852 69860 204916
rect 167316 204716 167380 204780
rect 231900 204716 231964 204780
rect 68324 203356 68388 203420
rect 69612 201180 69676 201244
rect 70164 200228 70228 200292
rect 67404 200092 67468 200156
rect 69244 200092 69308 200156
rect 68692 198732 68756 198796
rect 169892 198324 169956 198388
rect 119292 196692 119356 196756
rect 120212 196556 120276 196620
rect 167684 195196 167748 195260
rect 69796 194516 69860 194580
rect 167868 193156 167932 193220
rect 122236 192476 122300 192540
rect 69612 188940 69676 189004
rect 71268 180916 71332 180980
rect 71084 180780 71148 180844
rect 69244 179284 69308 179348
rect 71268 178060 71332 178124
rect 68508 177244 68572 177308
rect 69244 175884 69308 175948
rect 122420 175884 122484 175948
rect 169524 175476 169588 175540
rect 68324 173980 68388 174044
rect 169892 169492 169956 169556
rect 199332 168268 199396 168332
rect 120580 166968 120644 166972
rect 120580 166912 120630 166968
rect 120630 166912 120644 166968
rect 120580 166908 120644 166912
rect 119108 165548 119172 165612
rect 119660 125428 119724 125492
rect 118924 125292 118988 125356
rect 199516 124204 199580 124268
rect 121868 123388 121932 123452
rect 122052 122844 122116 122908
rect 170076 120668 170140 120732
rect 169892 120396 169956 120460
rect 169708 120124 169772 120188
rect 166028 119308 166092 119372
rect 200068 119368 200132 119372
rect 200068 119312 200118 119368
rect 200118 119312 200132 119368
rect 200068 119308 200132 119312
rect 199700 119036 199764 119100
rect 166948 118764 167012 118828
rect 200068 118628 200132 118692
rect 199700 118356 199764 118420
rect 166028 117948 166092 118012
rect 200068 117948 200132 118012
rect 199700 117676 199764 117740
rect 68876 117328 68940 117332
rect 68876 117272 68890 117328
rect 68890 117272 68940 117328
rect 68876 117268 68940 117272
rect 200068 117268 200132 117332
rect 199700 116996 199764 117060
rect 170260 116860 170324 116924
rect 166948 116452 167012 116516
rect 199516 116316 199580 116380
rect 200068 115908 200132 115972
rect 199700 115636 199764 115700
rect 200068 115228 200132 115292
rect 199700 114956 199764 115020
rect 170260 114820 170324 114884
rect 200068 114548 200132 114612
rect 170076 114004 170140 114068
rect 169892 113868 169956 113932
rect 169708 113732 169772 113796
rect 199700 113596 199764 113660
rect 200068 113188 200132 113252
rect 199700 112780 199764 112844
rect 70532 112508 70596 112572
rect 67220 112372 67284 112436
rect 200068 112508 200132 112572
rect 167500 112236 167564 112300
rect 199700 112100 199764 112164
rect 69428 111964 69492 112028
rect 70164 111828 70228 111892
rect 167316 111828 167380 111892
rect 200068 111828 200132 111892
rect 199700 111420 199764 111484
rect 70164 111284 70228 111348
rect 69060 110876 69124 110940
rect 106044 111148 106108 111212
rect 200068 111148 200132 111212
rect 105676 110876 105740 110940
rect 169340 110740 169404 110804
rect 199700 110740 199764 110804
rect 200068 110468 200132 110532
rect 106044 110332 106108 110396
rect 105676 110196 105740 110260
rect 199700 110060 199764 110124
rect 106044 109788 106108 109852
rect 200068 109788 200132 109852
rect 105676 109516 105740 109580
rect 199700 109380 199764 109444
rect 200068 109108 200132 109172
rect 106044 108972 106108 109036
rect 70348 108836 70412 108900
rect 105676 108836 105740 108900
rect 169892 108836 169956 108900
rect 106044 108428 106108 108492
rect 200068 108428 200132 108492
rect 105676 108156 105740 108220
rect 199700 108156 199764 108220
rect 105676 107340 105740 107404
rect 199700 107340 199764 107404
rect 106044 107068 106108 107132
rect 200068 107068 200132 107132
rect 105676 106660 105740 106724
rect 199700 106660 199764 106724
rect 106044 106388 106108 106452
rect 200068 106388 200132 106452
rect 105676 105980 105740 106044
rect 199516 105980 199580 106044
rect 106044 105708 106108 105772
rect 200068 105708 200132 105772
rect 199700 105436 199764 105500
rect 200068 105028 200132 105092
rect 105676 104756 105740 104820
rect 106044 104756 106108 104820
rect 199516 104620 199580 104684
rect 106044 104348 106108 104412
rect 200068 104408 200132 104412
rect 200068 104352 200118 104408
rect 200118 104352 200132 104408
rect 200068 104348 200132 104352
rect 105676 104076 105740 104140
rect 199700 104076 199764 104140
rect 200068 103668 200132 103732
rect 105676 103260 105740 103324
rect 106044 102988 106108 103052
rect 200068 102988 200132 103052
rect 199700 102716 199764 102780
rect 105676 102580 105740 102644
rect 106044 102308 106108 102372
rect 67220 102036 67284 102100
rect 105676 101900 105740 101964
rect 199700 101900 199764 101964
rect 106044 101628 106108 101692
rect 200068 101628 200132 101692
rect 105676 101220 105740 101284
rect 167500 101220 167564 101284
rect 169524 101220 169588 101284
rect 199700 101220 199764 101284
rect 106044 100948 106108 101012
rect 200068 100948 200132 101012
rect 201540 100948 201604 101012
rect 105676 100540 105740 100604
rect 199700 100540 199764 100604
rect 106044 100268 106108 100332
rect 200068 100268 200132 100332
rect 105676 99860 105740 99924
rect 199700 99860 199764 99924
rect 106044 99588 106108 99652
rect 200068 99588 200132 99652
rect 105676 99180 105740 99244
rect 106044 98908 106108 98972
rect 170076 98908 170140 98972
rect 199700 99180 199764 99244
rect 200068 98908 200132 98972
rect 199700 98500 199764 98564
rect 200068 98288 200132 98292
rect 200068 98232 200118 98288
rect 200118 98232 200132 98288
rect 200068 98228 200132 98232
rect 105676 97820 105740 97884
rect 106044 97820 106108 97884
rect 106044 97548 106108 97612
rect 200068 97548 200132 97612
rect 105492 97276 105556 97340
rect 199700 97276 199764 97340
rect 200068 96868 200132 96932
rect 105676 96596 105740 96660
rect 199700 96596 199764 96660
rect 106044 96460 106108 96524
rect 167500 96460 167564 96524
rect 106044 96188 106108 96252
rect 200068 96188 200132 96252
rect 105676 95916 105740 95980
rect 199700 95916 199764 95980
rect 167316 95780 167380 95844
rect 106044 95508 106108 95572
rect 200068 95508 200132 95572
rect 105676 95236 105740 95300
rect 120028 95296 120092 95300
rect 120028 95240 120042 95296
rect 120042 95240 120092 95296
rect 120028 95236 120092 95240
rect 199700 95236 199764 95300
rect 106044 94828 106108 94892
rect 200068 94828 200132 94892
rect 199700 94556 199764 94620
rect 105676 94420 105740 94484
rect 106044 94148 106108 94212
rect 200068 94148 200132 94212
rect 105492 93876 105556 93940
rect 199700 93876 199764 93940
rect 106044 93468 106108 93532
rect 105676 93196 105740 93260
rect 199700 93060 199764 93124
rect 106044 92788 106108 92852
rect 200068 92788 200132 92852
rect 69428 92516 69492 92580
rect 105676 92516 105740 92580
rect 200068 92108 200132 92172
rect 199700 91836 199764 91900
rect 106044 91428 106108 91492
rect 200068 91428 200132 91492
rect 201724 91428 201788 91492
rect 105676 91156 105740 91220
rect 199700 91156 199764 91220
rect 106044 90748 106108 90812
rect 200068 90748 200132 90812
rect 105676 90476 105740 90540
rect 199700 90476 199764 90540
rect 106044 90068 106108 90132
rect 200068 90068 200132 90132
rect 105676 89796 105740 89860
rect 199700 89796 199764 89860
rect 106044 89388 106108 89452
rect 200068 89388 200132 89452
rect 105676 89116 105740 89180
rect 199700 89116 199764 89180
rect 106044 88708 106108 88772
rect 200068 88708 200132 88772
rect 105676 88436 105740 88500
rect 199700 88436 199764 88500
rect 106044 88028 106108 88092
rect 200068 88028 200132 88092
rect 105676 87756 105740 87820
rect 199700 87756 199764 87820
rect 167684 87484 167748 87548
rect 106044 87348 106108 87412
rect 105676 87076 105740 87140
rect 106044 86668 106108 86732
rect 200068 86668 200132 86732
rect 105676 86396 105740 86460
rect 199700 86396 199764 86460
rect 106044 85988 106108 86052
rect 200068 86048 200132 86052
rect 200068 85992 200118 86048
rect 200118 85992 200132 86048
rect 200068 85988 200132 85992
rect 105676 85716 105740 85780
rect 199700 85580 199764 85644
rect 200068 85640 200132 85644
rect 200068 85584 200118 85640
rect 200118 85584 200132 85640
rect 200068 85580 200132 85584
rect 167868 85036 167932 85100
rect 69060 84900 69124 84964
rect 199700 84900 199764 84964
rect 200068 84764 200132 84828
rect 106044 84628 106108 84692
rect 105676 84356 105740 84420
rect 199700 84220 199764 84284
rect 200068 84220 200132 84284
rect 106044 83948 106108 84012
rect 105676 83676 105740 83740
rect 68692 83540 68756 83604
rect 106044 83268 106108 83332
rect 199332 83540 199396 83604
rect 106780 83132 106844 83196
rect 200068 83268 200132 83332
rect 105676 82996 105740 83060
rect 199700 82996 199764 83060
rect 200068 82860 200132 82924
rect 106044 82588 106108 82652
rect 105676 82316 105740 82380
rect 106044 81908 106108 81972
rect 199700 82180 199764 82244
rect 106228 81772 106292 81836
rect 200068 81908 200132 81972
rect 105676 81636 105740 81700
rect 106044 81228 106108 81292
rect 105676 80956 105740 81020
rect 199700 80820 199764 80884
rect 106044 80548 106108 80612
rect 200068 80548 200132 80612
rect 105676 80276 105740 80340
rect 199700 80140 199764 80204
rect 200068 80004 200132 80068
rect 106044 79868 106108 79932
rect 105676 79596 105740 79660
rect 199700 79460 199764 79524
rect 106044 79188 106108 79252
rect 200068 79188 200132 79252
rect 105676 78916 105740 78980
rect 199700 78780 199764 78844
rect 200068 78644 200132 78708
rect 199332 78100 199396 78164
rect 106044 77828 106108 77892
rect 105676 77556 105740 77620
rect 199700 77420 199764 77484
rect 200068 77284 200132 77348
rect 105676 76740 105740 76804
rect 199700 76740 199764 76804
rect 106044 76468 106108 76532
rect 106412 76468 106476 76532
rect 200068 76468 200132 76532
rect 105676 76060 105740 76124
rect 106044 75924 106108 75988
rect 67404 75652 67468 75716
rect 68876 75652 68940 75716
rect 106044 75652 106108 75716
rect 105676 75516 105740 75580
rect 199700 75380 199764 75444
rect 106044 75108 106108 75172
rect 200068 75108 200132 75172
rect 106228 75032 106292 75036
rect 106228 74976 106242 75032
rect 106242 74976 106292 75032
rect 106228 74972 106292 74976
rect 105676 74836 105740 74900
rect 199332 74700 199396 74764
rect 200068 74700 200132 74764
rect 68508 74020 68572 74084
rect 105676 74020 105740 74084
rect 106044 74020 106108 74084
rect 199700 74020 199764 74084
rect 168972 73884 169036 73948
rect 170260 73748 170324 73812
rect 200068 73748 200132 73812
rect 106044 73612 106108 73676
rect 69244 73340 69308 73404
rect 68324 73204 68388 73268
rect 105676 73340 105740 73404
rect 199700 73340 199764 73404
rect 70532 73204 70596 73268
rect 200068 73204 200132 73268
rect 106044 72796 106108 72860
rect 105676 72660 105740 72724
rect 167868 72660 167932 72724
rect 199700 72660 199764 72724
rect 200068 72388 200132 72452
rect 106044 72252 106108 72316
rect 105676 72116 105740 72180
rect 199700 71980 199764 72044
rect 200068 71844 200132 71908
rect 106044 71028 106108 71092
rect 105676 70620 105740 70684
rect 106044 70212 106108 70276
rect 105676 70076 105740 70140
rect 70532 69940 70596 70004
rect 69060 69804 69124 69868
rect 167684 69804 167748 69868
rect 168972 69804 169036 69868
rect 167316 69668 167380 69732
rect 170260 69668 170324 69732
rect 68692 69532 68756 69596
rect 106780 69532 106844 69596
rect 201724 69532 201788 69596
rect 68876 69396 68940 69460
rect 106044 69396 106108 69460
rect 199332 69396 199396 69460
rect 105492 69260 105556 69324
rect 199148 69260 199212 69324
rect 200068 68852 200132 68916
rect 105308 67220 105372 67284
rect 201540 67220 201604 67284
rect 167868 64772 167932 64836
rect 167868 58516 167932 58580
rect 170076 57156 170140 57220
rect 167500 54436 167564 54500
rect 169340 53076 169404 53140
rect 169708 43420 169772 43484
rect 169892 40564 169956 40628
rect 169524 19892 169588 19956
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 677494 -8106 711002
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 -8106 677494
rect -8726 677174 -8106 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 -8106 677174
rect -8726 641494 -8106 676938
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 -8106 641494
rect -8726 641174 -8106 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 -8106 641174
rect -8726 605494 -8106 640938
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 -8106 605494
rect -8726 605174 -8106 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 -8106 605174
rect -8726 569494 -8106 604938
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 -8106 569494
rect -8726 569174 -8106 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 -8106 569174
rect -8726 533494 -8106 568938
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 -8106 533494
rect -8726 533174 -8106 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 -8106 533174
rect -8726 497494 -8106 532938
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 -8106 497494
rect -8726 497174 -8106 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 -8106 497174
rect -8726 461494 -8106 496938
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 -8106 461494
rect -8726 461174 -8106 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 -8106 461174
rect -8726 425494 -8106 460938
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 -8106 425494
rect -8726 425174 -8106 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 -8106 425174
rect -8726 389494 -8106 424938
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 -8106 389494
rect -8726 389174 -8106 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 -8106 389174
rect -8726 353494 -8106 388938
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 -8106 353494
rect -8726 353174 -8106 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 -8106 353174
rect -8726 317494 -8106 352938
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 -8106 317494
rect -8726 317174 -8106 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 -8106 317174
rect -8726 281494 -8106 316938
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 -8106 281494
rect -8726 281174 -8106 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 -8106 281174
rect -8726 245494 -8106 280938
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 -8106 245494
rect -8726 245174 -8106 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 -8106 245174
rect -8726 209494 -8106 244938
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 -8106 209494
rect -8726 209174 -8106 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 -8106 209174
rect -8726 173494 -8106 208938
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 -8106 173494
rect -8726 173174 -8106 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 -8106 173174
rect -8726 137494 -8106 172938
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 -8106 137494
rect -8726 137174 -8106 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 -8106 137174
rect -8726 101494 -8106 136938
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 -8106 101494
rect -8726 101174 -8106 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 -8106 101174
rect -8726 65494 -8106 100938
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 -8106 65494
rect -8726 65174 -8106 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 -8106 65174
rect -8726 29494 -8106 64938
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 -8106 29494
rect -8726 29174 -8106 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 -8106 29174
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 673774 -7146 710042
rect -7766 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 -7146 673774
rect -7766 673454 -7146 673538
rect -7766 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 -7146 673454
rect -7766 637774 -7146 673218
rect -7766 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 -7146 637774
rect -7766 637454 -7146 637538
rect -7766 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 -7146 637454
rect -7766 601774 -7146 637218
rect -7766 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 -7146 601774
rect -7766 601454 -7146 601538
rect -7766 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 -7146 601454
rect -7766 565774 -7146 601218
rect -7766 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 -7146 565774
rect -7766 565454 -7146 565538
rect -7766 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 -7146 565454
rect -7766 529774 -7146 565218
rect -7766 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 -7146 529774
rect -7766 529454 -7146 529538
rect -7766 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 -7146 529454
rect -7766 493774 -7146 529218
rect -7766 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 -7146 493774
rect -7766 493454 -7146 493538
rect -7766 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 -7146 493454
rect -7766 457774 -7146 493218
rect -7766 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 -7146 457774
rect -7766 457454 -7146 457538
rect -7766 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 -7146 457454
rect -7766 421774 -7146 457218
rect -7766 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 -7146 421774
rect -7766 421454 -7146 421538
rect -7766 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 -7146 421454
rect -7766 385774 -7146 421218
rect -7766 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 -7146 385774
rect -7766 385454 -7146 385538
rect -7766 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 -7146 385454
rect -7766 349774 -7146 385218
rect -7766 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 -7146 349774
rect -7766 349454 -7146 349538
rect -7766 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 -7146 349454
rect -7766 313774 -7146 349218
rect -7766 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 -7146 313774
rect -7766 313454 -7146 313538
rect -7766 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 -7146 313454
rect -7766 277774 -7146 313218
rect -7766 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 -7146 277774
rect -7766 277454 -7146 277538
rect -7766 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 -7146 277454
rect -7766 241774 -7146 277218
rect -7766 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 -7146 241774
rect -7766 241454 -7146 241538
rect -7766 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 -7146 241454
rect -7766 205774 -7146 241218
rect -7766 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 -7146 205774
rect -7766 205454 -7146 205538
rect -7766 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 -7146 205454
rect -7766 169774 -7146 205218
rect -7766 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 -7146 169774
rect -7766 169454 -7146 169538
rect -7766 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 -7146 169454
rect -7766 133774 -7146 169218
rect -7766 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 -7146 133774
rect -7766 133454 -7146 133538
rect -7766 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 -7146 133454
rect -7766 97774 -7146 133218
rect -7766 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 -7146 97774
rect -7766 97454 -7146 97538
rect -7766 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 -7146 97454
rect -7766 61774 -7146 97218
rect -7766 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 -7146 61774
rect -7766 61454 -7146 61538
rect -7766 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 -7146 61454
rect -7766 25774 -7146 61218
rect -7766 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 -7146 25774
rect -7766 25454 -7146 25538
rect -7766 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 -7146 25454
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 670054 -6186 709082
rect -6806 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 -6186 670054
rect -6806 669734 -6186 669818
rect -6806 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 -6186 669734
rect -6806 634054 -6186 669498
rect -6806 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 -6186 634054
rect -6806 633734 -6186 633818
rect -6806 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 -6186 633734
rect -6806 598054 -6186 633498
rect -6806 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 -6186 598054
rect -6806 597734 -6186 597818
rect -6806 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 -6186 597734
rect -6806 562054 -6186 597498
rect -6806 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 -6186 562054
rect -6806 561734 -6186 561818
rect -6806 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 -6186 561734
rect -6806 526054 -6186 561498
rect -6806 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 -6186 526054
rect -6806 525734 -6186 525818
rect -6806 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 -6186 525734
rect -6806 490054 -6186 525498
rect -6806 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 -6186 490054
rect -6806 489734 -6186 489818
rect -6806 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 -6186 489734
rect -6806 454054 -6186 489498
rect -6806 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 -6186 454054
rect -6806 453734 -6186 453818
rect -6806 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 -6186 453734
rect -6806 418054 -6186 453498
rect -6806 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 -6186 418054
rect -6806 417734 -6186 417818
rect -6806 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 -6186 417734
rect -6806 382054 -6186 417498
rect -6806 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 -6186 382054
rect -6806 381734 -6186 381818
rect -6806 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 -6186 381734
rect -6806 346054 -6186 381498
rect -6806 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 -6186 346054
rect -6806 345734 -6186 345818
rect -6806 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 -6186 345734
rect -6806 310054 -6186 345498
rect -6806 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 -6186 310054
rect -6806 309734 -6186 309818
rect -6806 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 -6186 309734
rect -6806 274054 -6186 309498
rect -6806 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 -6186 274054
rect -6806 273734 -6186 273818
rect -6806 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 -6186 273734
rect -6806 238054 -6186 273498
rect -6806 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 -6186 238054
rect -6806 237734 -6186 237818
rect -6806 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 -6186 237734
rect -6806 202054 -6186 237498
rect -6806 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 -6186 202054
rect -6806 201734 -6186 201818
rect -6806 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 -6186 201734
rect -6806 166054 -6186 201498
rect -6806 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 -6186 166054
rect -6806 165734 -6186 165818
rect -6806 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 -6186 165734
rect -6806 130054 -6186 165498
rect -6806 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 -6186 130054
rect -6806 129734 -6186 129818
rect -6806 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 -6186 129734
rect -6806 94054 -6186 129498
rect -6806 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 -6186 94054
rect -6806 93734 -6186 93818
rect -6806 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 -6186 93734
rect -6806 58054 -6186 93498
rect -6806 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 -6186 58054
rect -6806 57734 -6186 57818
rect -6806 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 -6186 57734
rect -6806 22054 -6186 57498
rect -6806 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 -6186 22054
rect -6806 21734 -6186 21818
rect -6806 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 -6186 21734
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 666334 -5226 708122
rect -5846 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 -5226 666334
rect -5846 666014 -5226 666098
rect -5846 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 -5226 666014
rect -5846 630334 -5226 665778
rect -5846 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 -5226 630334
rect -5846 630014 -5226 630098
rect -5846 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 -5226 630014
rect -5846 594334 -5226 629778
rect -5846 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 -5226 594334
rect -5846 594014 -5226 594098
rect -5846 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 -5226 594014
rect -5846 558334 -5226 593778
rect -5846 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 -5226 558334
rect -5846 558014 -5226 558098
rect -5846 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 -5226 558014
rect -5846 522334 -5226 557778
rect -5846 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 -5226 522334
rect -5846 522014 -5226 522098
rect -5846 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 -5226 522014
rect -5846 486334 -5226 521778
rect -5846 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 -5226 486334
rect -5846 486014 -5226 486098
rect -5846 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 -5226 486014
rect -5846 450334 -5226 485778
rect -5846 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 -5226 450334
rect -5846 450014 -5226 450098
rect -5846 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 -5226 450014
rect -5846 414334 -5226 449778
rect -5846 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 -5226 414334
rect -5846 414014 -5226 414098
rect -5846 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 -5226 414014
rect -5846 378334 -5226 413778
rect -5846 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 -5226 378334
rect -5846 378014 -5226 378098
rect -5846 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 -5226 378014
rect -5846 342334 -5226 377778
rect -5846 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 -5226 342334
rect -5846 342014 -5226 342098
rect -5846 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 -5226 342014
rect -5846 306334 -5226 341778
rect -5846 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 -5226 306334
rect -5846 306014 -5226 306098
rect -5846 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 -5226 306014
rect -5846 270334 -5226 305778
rect -5846 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 -5226 270334
rect -5846 270014 -5226 270098
rect -5846 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 -5226 270014
rect -5846 234334 -5226 269778
rect -5846 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 -5226 234334
rect -5846 234014 -5226 234098
rect -5846 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 -5226 234014
rect -5846 198334 -5226 233778
rect -5846 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 -5226 198334
rect -5846 198014 -5226 198098
rect -5846 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 -5226 198014
rect -5846 162334 -5226 197778
rect -5846 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 -5226 162334
rect -5846 162014 -5226 162098
rect -5846 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 -5226 162014
rect -5846 126334 -5226 161778
rect -5846 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 -5226 126334
rect -5846 126014 -5226 126098
rect -5846 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 -5226 126014
rect -5846 90334 -5226 125778
rect -5846 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 -5226 90334
rect -5846 90014 -5226 90098
rect -5846 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 -5226 90014
rect -5846 54334 -5226 89778
rect -5846 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 -5226 54334
rect -5846 54014 -5226 54098
rect -5846 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 -5226 54014
rect -5846 18334 -5226 53778
rect -5846 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 -5226 18334
rect -5846 18014 -5226 18098
rect -5846 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 -5226 18014
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 698614 -4266 707162
rect -4886 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 -4266 698614
rect -4886 698294 -4266 698378
rect -4886 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 -4266 698294
rect -4886 662614 -4266 698058
rect -4886 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 -4266 662614
rect -4886 662294 -4266 662378
rect -4886 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 -4266 662294
rect -4886 626614 -4266 662058
rect -4886 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 -4266 626614
rect -4886 626294 -4266 626378
rect -4886 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 -4266 626294
rect -4886 590614 -4266 626058
rect -4886 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 -4266 590614
rect -4886 590294 -4266 590378
rect -4886 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 -4266 590294
rect -4886 554614 -4266 590058
rect -4886 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 -4266 554614
rect -4886 554294 -4266 554378
rect -4886 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 -4266 554294
rect -4886 518614 -4266 554058
rect -4886 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 -4266 518614
rect -4886 518294 -4266 518378
rect -4886 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 -4266 518294
rect -4886 482614 -4266 518058
rect -4886 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 -4266 482614
rect -4886 482294 -4266 482378
rect -4886 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 -4266 482294
rect -4886 446614 -4266 482058
rect -4886 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 -4266 446614
rect -4886 446294 -4266 446378
rect -4886 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 -4266 446294
rect -4886 410614 -4266 446058
rect -4886 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 -4266 410614
rect -4886 410294 -4266 410378
rect -4886 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 -4266 410294
rect -4886 374614 -4266 410058
rect -4886 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 -4266 374614
rect -4886 374294 -4266 374378
rect -4886 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 -4266 374294
rect -4886 338614 -4266 374058
rect -4886 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 -4266 338614
rect -4886 338294 -4266 338378
rect -4886 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 -4266 338294
rect -4886 302614 -4266 338058
rect -4886 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 -4266 302614
rect -4886 302294 -4266 302378
rect -4886 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 -4266 302294
rect -4886 266614 -4266 302058
rect -4886 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 -4266 266614
rect -4886 266294 -4266 266378
rect -4886 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 -4266 266294
rect -4886 230614 -4266 266058
rect -4886 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 -4266 230614
rect -4886 230294 -4266 230378
rect -4886 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 -4266 230294
rect -4886 194614 -4266 230058
rect -4886 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 -4266 194614
rect -4886 194294 -4266 194378
rect -4886 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 -4266 194294
rect -4886 158614 -4266 194058
rect -4886 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 -4266 158614
rect -4886 158294 -4266 158378
rect -4886 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 -4266 158294
rect -4886 122614 -4266 158058
rect -4886 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 -4266 122614
rect -4886 122294 -4266 122378
rect -4886 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 -4266 122294
rect -4886 86614 -4266 122058
rect -4886 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 -4266 86614
rect -4886 86294 -4266 86378
rect -4886 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 -4266 86294
rect -4886 50614 -4266 86058
rect -4886 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 -4266 50614
rect -4886 50294 -4266 50378
rect -4886 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 -4266 50294
rect -4886 14614 -4266 50058
rect -4886 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 -4266 14614
rect -4886 14294 -4266 14378
rect -4886 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 -4266 14294
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 694894 -3306 706202
rect -3926 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 -3306 694894
rect -3926 694574 -3306 694658
rect -3926 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 -3306 694574
rect -3926 658894 -3306 694338
rect -3926 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 -3306 658894
rect -3926 658574 -3306 658658
rect -3926 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 -3306 658574
rect -3926 622894 -3306 658338
rect -3926 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 -3306 622894
rect -3926 622574 -3306 622658
rect -3926 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 -3306 622574
rect -3926 586894 -3306 622338
rect -3926 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 -3306 586894
rect -3926 586574 -3306 586658
rect -3926 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 -3306 586574
rect -3926 550894 -3306 586338
rect -3926 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 -3306 550894
rect -3926 550574 -3306 550658
rect -3926 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 -3306 550574
rect -3926 514894 -3306 550338
rect -3926 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 -3306 514894
rect -3926 514574 -3306 514658
rect -3926 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 -3306 514574
rect -3926 478894 -3306 514338
rect -3926 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 -3306 478894
rect -3926 478574 -3306 478658
rect -3926 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 -3306 478574
rect -3926 442894 -3306 478338
rect -3926 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 -3306 442894
rect -3926 442574 -3306 442658
rect -3926 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 -3306 442574
rect -3926 406894 -3306 442338
rect -3926 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 -3306 406894
rect -3926 406574 -3306 406658
rect -3926 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 -3306 406574
rect -3926 370894 -3306 406338
rect -3926 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 -3306 370894
rect -3926 370574 -3306 370658
rect -3926 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 -3306 370574
rect -3926 334894 -3306 370338
rect -3926 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 -3306 334894
rect -3926 334574 -3306 334658
rect -3926 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 -3306 334574
rect -3926 298894 -3306 334338
rect -3926 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 -3306 298894
rect -3926 298574 -3306 298658
rect -3926 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 -3306 298574
rect -3926 262894 -3306 298338
rect -3926 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 -3306 262894
rect -3926 262574 -3306 262658
rect -3926 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 -3306 262574
rect -3926 226894 -3306 262338
rect -3926 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 -3306 226894
rect -3926 226574 -3306 226658
rect -3926 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 -3306 226574
rect -3926 190894 -3306 226338
rect -3926 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 -3306 190894
rect -3926 190574 -3306 190658
rect -3926 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 -3306 190574
rect -3926 154894 -3306 190338
rect -3926 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 -3306 154894
rect -3926 154574 -3306 154658
rect -3926 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 -3306 154574
rect -3926 118894 -3306 154338
rect -3926 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 -3306 118894
rect -3926 118574 -3306 118658
rect -3926 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 -3306 118574
rect -3926 82894 -3306 118338
rect -3926 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 -3306 82894
rect -3926 82574 -3306 82658
rect -3926 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 -3306 82574
rect -3926 46894 -3306 82338
rect -3926 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 -3306 46894
rect -3926 46574 -3306 46658
rect -3926 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 -3306 46574
rect -3926 10894 -3306 46338
rect -3926 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 -3306 10894
rect -3926 10574 -3306 10658
rect -3926 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 -3306 10574
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691174 -2346 705242
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 -2346 691174
rect -2966 690854 -2346 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 -2346 690854
rect -2966 655174 -2346 690618
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 -2346 655174
rect -2966 654854 -2346 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 -2346 654854
rect -2966 619174 -2346 654618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 583174 -2346 618618
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 -2346 583174
rect -2966 582854 -2346 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 -2346 582854
rect -2966 547174 -2346 582618
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 -2346 547174
rect -2966 546854 -2346 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 -2346 546854
rect -2966 511174 -2346 546618
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 -2346 511174
rect -2966 510854 -2346 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 -2346 510854
rect -2966 475174 -2346 510618
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 -2346 475174
rect -2966 474854 -2346 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 -2346 474854
rect -2966 439174 -2346 474618
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 -2346 439174
rect -2966 438854 -2346 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 -2346 438854
rect -2966 403174 -2346 438618
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 -2346 403174
rect -2966 402854 -2346 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 -2346 402854
rect -2966 367174 -2346 402618
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 -2346 367174
rect -2966 366854 -2346 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 -2346 366854
rect -2966 331174 -2346 366618
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 -2346 331174
rect -2966 330854 -2346 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 -2346 330854
rect -2966 295174 -2346 330618
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 -2346 295174
rect -2966 294854 -2346 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 -2346 294854
rect -2966 259174 -2346 294618
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 -2346 259174
rect -2966 258854 -2346 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 -2346 258854
rect -2966 223174 -2346 258618
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 -2346 223174
rect -2966 222854 -2346 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 -2346 222854
rect -2966 187174 -2346 222618
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 -2346 187174
rect -2966 186854 -2346 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 -2346 186854
rect -2966 151174 -2346 186618
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 -2346 151174
rect -2966 150854 -2346 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 -2346 150854
rect -2966 115174 -2346 150618
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 -2346 115174
rect -2966 114854 -2346 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 -2346 114854
rect -2966 79174 -2346 114618
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 -2346 79174
rect -2966 78854 -2346 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 -2346 78854
rect -2966 43174 -2346 78618
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 -2346 43174
rect -2966 42854 -2346 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 -2346 42854
rect -2966 7174 -2346 42618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 705798 6134 711590
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 691174 6134 705242
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 5514 -1306 6134 6618
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -7654 6134 -1862
rect 9234 706758 9854 711590
rect 9234 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 9854 706758
rect 9234 706438 9854 706522
rect 9234 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 9854 706438
rect 9234 694894 9854 706202
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect 9234 -2266 9854 10338
rect 9234 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 9854 -2266
rect 9234 -2586 9854 -2502
rect 9234 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 9854 -2586
rect 9234 -7654 9854 -2822
rect 12954 707718 13574 711590
rect 12954 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 13574 707718
rect 12954 707398 13574 707482
rect 12954 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 13574 707398
rect 12954 698614 13574 707162
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect 12954 -3226 13574 14058
rect 12954 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 13574 -3226
rect 12954 -3546 13574 -3462
rect 12954 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 13574 -3546
rect 12954 -7654 13574 -3782
rect 16674 708678 17294 711590
rect 16674 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 17294 708678
rect 16674 708358 17294 708442
rect 16674 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 17294 708358
rect 16674 666334 17294 708122
rect 16674 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 17294 666334
rect 16674 666014 17294 666098
rect 16674 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 17294 666014
rect 16674 630334 17294 665778
rect 16674 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 17294 630334
rect 16674 630014 17294 630098
rect 16674 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 17294 630014
rect 16674 594334 17294 629778
rect 16674 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 17294 594334
rect 16674 594014 17294 594098
rect 16674 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 17294 594014
rect 16674 558334 17294 593778
rect 16674 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 17294 558334
rect 16674 558014 17294 558098
rect 16674 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 17294 558014
rect 16674 522334 17294 557778
rect 16674 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 17294 522334
rect 16674 522014 17294 522098
rect 16674 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 17294 522014
rect 16674 486334 17294 521778
rect 16674 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 17294 486334
rect 16674 486014 17294 486098
rect 16674 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 17294 486014
rect 16674 450334 17294 485778
rect 16674 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 17294 450334
rect 16674 450014 17294 450098
rect 16674 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 17294 450014
rect 16674 414334 17294 449778
rect 16674 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 17294 414334
rect 16674 414014 17294 414098
rect 16674 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 17294 414014
rect 16674 378334 17294 413778
rect 16674 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 17294 378334
rect 16674 378014 17294 378098
rect 16674 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 17294 378014
rect 16674 342334 17294 377778
rect 16674 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 17294 342334
rect 16674 342014 17294 342098
rect 16674 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 17294 342014
rect 16674 306334 17294 341778
rect 16674 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 17294 306334
rect 16674 306014 17294 306098
rect 16674 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 17294 306014
rect 16674 270334 17294 305778
rect 16674 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 17294 270334
rect 16674 270014 17294 270098
rect 16674 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 17294 270014
rect 16674 234334 17294 269778
rect 16674 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 17294 234334
rect 16674 234014 17294 234098
rect 16674 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 17294 234014
rect 16674 198334 17294 233778
rect 16674 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 17294 198334
rect 16674 198014 17294 198098
rect 16674 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 17294 198014
rect 16674 162334 17294 197778
rect 16674 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 17294 162334
rect 16674 162014 17294 162098
rect 16674 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 17294 162014
rect 16674 126334 17294 161778
rect 16674 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 17294 126334
rect 16674 126014 17294 126098
rect 16674 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 17294 126014
rect 16674 90334 17294 125778
rect 16674 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 17294 90334
rect 16674 90014 17294 90098
rect 16674 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 17294 90014
rect 16674 54334 17294 89778
rect 16674 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 17294 54334
rect 16674 54014 17294 54098
rect 16674 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 17294 54014
rect 16674 18334 17294 53778
rect 16674 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 17294 18334
rect 16674 18014 17294 18098
rect 16674 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 17294 18014
rect 16674 -4186 17294 17778
rect 16674 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 17294 -4186
rect 16674 -4506 17294 -4422
rect 16674 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 17294 -4506
rect 16674 -7654 17294 -4742
rect 20394 709638 21014 711590
rect 20394 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 21014 709638
rect 20394 709318 21014 709402
rect 20394 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 21014 709318
rect 20394 670054 21014 709082
rect 20394 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 21014 670054
rect 20394 669734 21014 669818
rect 20394 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 21014 669734
rect 20394 634054 21014 669498
rect 20394 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 21014 634054
rect 20394 633734 21014 633818
rect 20394 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 21014 633734
rect 20394 598054 21014 633498
rect 20394 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 21014 598054
rect 20394 597734 21014 597818
rect 20394 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 21014 597734
rect 20394 562054 21014 597498
rect 20394 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 21014 562054
rect 20394 561734 21014 561818
rect 20394 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 21014 561734
rect 20394 526054 21014 561498
rect 20394 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 21014 526054
rect 20394 525734 21014 525818
rect 20394 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 21014 525734
rect 20394 490054 21014 525498
rect 20394 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 21014 490054
rect 20394 489734 21014 489818
rect 20394 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 21014 489734
rect 20394 454054 21014 489498
rect 20394 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 21014 454054
rect 20394 453734 21014 453818
rect 20394 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 21014 453734
rect 20394 418054 21014 453498
rect 20394 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 21014 418054
rect 20394 417734 21014 417818
rect 20394 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 21014 417734
rect 20394 382054 21014 417498
rect 20394 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 21014 382054
rect 20394 381734 21014 381818
rect 20394 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 21014 381734
rect 20394 346054 21014 381498
rect 20394 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 21014 346054
rect 20394 345734 21014 345818
rect 20394 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 21014 345734
rect 20394 310054 21014 345498
rect 20394 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 21014 310054
rect 20394 309734 21014 309818
rect 20394 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 21014 309734
rect 20394 274054 21014 309498
rect 20394 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 21014 274054
rect 20394 273734 21014 273818
rect 20394 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 21014 273734
rect 20394 238054 21014 273498
rect 20394 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 21014 238054
rect 20394 237734 21014 237818
rect 20394 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 21014 237734
rect 20394 202054 21014 237498
rect 20394 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 21014 202054
rect 20394 201734 21014 201818
rect 20394 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 21014 201734
rect 20394 166054 21014 201498
rect 20394 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 21014 166054
rect 20394 165734 21014 165818
rect 20394 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 21014 165734
rect 20394 130054 21014 165498
rect 20394 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 21014 130054
rect 20394 129734 21014 129818
rect 20394 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 21014 129734
rect 20394 94054 21014 129498
rect 20394 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 21014 94054
rect 20394 93734 21014 93818
rect 20394 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 21014 93734
rect 20394 58054 21014 93498
rect 20394 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 21014 58054
rect 20394 57734 21014 57818
rect 20394 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 21014 57734
rect 20394 22054 21014 57498
rect 20394 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 21014 22054
rect 20394 21734 21014 21818
rect 20394 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 21014 21734
rect 20394 -5146 21014 21498
rect 20394 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 21014 -5146
rect 20394 -5466 21014 -5382
rect 20394 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 21014 -5466
rect 20394 -7654 21014 -5702
rect 24114 710598 24734 711590
rect 24114 710362 24146 710598
rect 24382 710362 24466 710598
rect 24702 710362 24734 710598
rect 24114 710278 24734 710362
rect 24114 710042 24146 710278
rect 24382 710042 24466 710278
rect 24702 710042 24734 710278
rect 24114 673774 24734 710042
rect 24114 673538 24146 673774
rect 24382 673538 24466 673774
rect 24702 673538 24734 673774
rect 24114 673454 24734 673538
rect 24114 673218 24146 673454
rect 24382 673218 24466 673454
rect 24702 673218 24734 673454
rect 24114 637774 24734 673218
rect 24114 637538 24146 637774
rect 24382 637538 24466 637774
rect 24702 637538 24734 637774
rect 24114 637454 24734 637538
rect 24114 637218 24146 637454
rect 24382 637218 24466 637454
rect 24702 637218 24734 637454
rect 24114 601774 24734 637218
rect 24114 601538 24146 601774
rect 24382 601538 24466 601774
rect 24702 601538 24734 601774
rect 24114 601454 24734 601538
rect 24114 601218 24146 601454
rect 24382 601218 24466 601454
rect 24702 601218 24734 601454
rect 24114 565774 24734 601218
rect 24114 565538 24146 565774
rect 24382 565538 24466 565774
rect 24702 565538 24734 565774
rect 24114 565454 24734 565538
rect 24114 565218 24146 565454
rect 24382 565218 24466 565454
rect 24702 565218 24734 565454
rect 24114 529774 24734 565218
rect 24114 529538 24146 529774
rect 24382 529538 24466 529774
rect 24702 529538 24734 529774
rect 24114 529454 24734 529538
rect 24114 529218 24146 529454
rect 24382 529218 24466 529454
rect 24702 529218 24734 529454
rect 24114 493774 24734 529218
rect 24114 493538 24146 493774
rect 24382 493538 24466 493774
rect 24702 493538 24734 493774
rect 24114 493454 24734 493538
rect 24114 493218 24146 493454
rect 24382 493218 24466 493454
rect 24702 493218 24734 493454
rect 24114 457774 24734 493218
rect 24114 457538 24146 457774
rect 24382 457538 24466 457774
rect 24702 457538 24734 457774
rect 24114 457454 24734 457538
rect 24114 457218 24146 457454
rect 24382 457218 24466 457454
rect 24702 457218 24734 457454
rect 24114 421774 24734 457218
rect 24114 421538 24146 421774
rect 24382 421538 24466 421774
rect 24702 421538 24734 421774
rect 24114 421454 24734 421538
rect 24114 421218 24146 421454
rect 24382 421218 24466 421454
rect 24702 421218 24734 421454
rect 24114 385774 24734 421218
rect 24114 385538 24146 385774
rect 24382 385538 24466 385774
rect 24702 385538 24734 385774
rect 24114 385454 24734 385538
rect 24114 385218 24146 385454
rect 24382 385218 24466 385454
rect 24702 385218 24734 385454
rect 24114 349774 24734 385218
rect 24114 349538 24146 349774
rect 24382 349538 24466 349774
rect 24702 349538 24734 349774
rect 24114 349454 24734 349538
rect 24114 349218 24146 349454
rect 24382 349218 24466 349454
rect 24702 349218 24734 349454
rect 24114 313774 24734 349218
rect 24114 313538 24146 313774
rect 24382 313538 24466 313774
rect 24702 313538 24734 313774
rect 24114 313454 24734 313538
rect 24114 313218 24146 313454
rect 24382 313218 24466 313454
rect 24702 313218 24734 313454
rect 24114 277774 24734 313218
rect 24114 277538 24146 277774
rect 24382 277538 24466 277774
rect 24702 277538 24734 277774
rect 24114 277454 24734 277538
rect 24114 277218 24146 277454
rect 24382 277218 24466 277454
rect 24702 277218 24734 277454
rect 24114 241774 24734 277218
rect 24114 241538 24146 241774
rect 24382 241538 24466 241774
rect 24702 241538 24734 241774
rect 24114 241454 24734 241538
rect 24114 241218 24146 241454
rect 24382 241218 24466 241454
rect 24702 241218 24734 241454
rect 24114 205774 24734 241218
rect 24114 205538 24146 205774
rect 24382 205538 24466 205774
rect 24702 205538 24734 205774
rect 24114 205454 24734 205538
rect 24114 205218 24146 205454
rect 24382 205218 24466 205454
rect 24702 205218 24734 205454
rect 24114 169774 24734 205218
rect 24114 169538 24146 169774
rect 24382 169538 24466 169774
rect 24702 169538 24734 169774
rect 24114 169454 24734 169538
rect 24114 169218 24146 169454
rect 24382 169218 24466 169454
rect 24702 169218 24734 169454
rect 24114 133774 24734 169218
rect 24114 133538 24146 133774
rect 24382 133538 24466 133774
rect 24702 133538 24734 133774
rect 24114 133454 24734 133538
rect 24114 133218 24146 133454
rect 24382 133218 24466 133454
rect 24702 133218 24734 133454
rect 24114 97774 24734 133218
rect 24114 97538 24146 97774
rect 24382 97538 24466 97774
rect 24702 97538 24734 97774
rect 24114 97454 24734 97538
rect 24114 97218 24146 97454
rect 24382 97218 24466 97454
rect 24702 97218 24734 97454
rect 24114 61774 24734 97218
rect 24114 61538 24146 61774
rect 24382 61538 24466 61774
rect 24702 61538 24734 61774
rect 24114 61454 24734 61538
rect 24114 61218 24146 61454
rect 24382 61218 24466 61454
rect 24702 61218 24734 61454
rect 24114 25774 24734 61218
rect 24114 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 24734 25774
rect 24114 25454 24734 25538
rect 24114 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 24734 25454
rect 24114 -6106 24734 25218
rect 24114 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 24734 -6106
rect 24114 -6426 24734 -6342
rect 24114 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 24734 -6426
rect 24114 -7654 24734 -6662
rect 27834 711558 28454 711590
rect 27834 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 28454 711558
rect 27834 711238 28454 711322
rect 27834 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 28454 711238
rect 27834 677494 28454 711002
rect 27834 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 28454 677494
rect 27834 677174 28454 677258
rect 27834 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 28454 677174
rect 27834 641494 28454 676938
rect 27834 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 28454 641494
rect 27834 641174 28454 641258
rect 27834 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 28454 641174
rect 27834 605494 28454 640938
rect 27834 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 28454 605494
rect 27834 605174 28454 605258
rect 27834 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 28454 605174
rect 27834 569494 28454 604938
rect 27834 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 28454 569494
rect 27834 569174 28454 569258
rect 27834 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 28454 569174
rect 27834 533494 28454 568938
rect 27834 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 28454 533494
rect 27834 533174 28454 533258
rect 27834 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 28454 533174
rect 27834 497494 28454 532938
rect 27834 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 28454 497494
rect 27834 497174 28454 497258
rect 27834 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 28454 497174
rect 27834 461494 28454 496938
rect 27834 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 28454 461494
rect 27834 461174 28454 461258
rect 27834 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 28454 461174
rect 27834 425494 28454 460938
rect 27834 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 28454 425494
rect 27834 425174 28454 425258
rect 27834 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 28454 425174
rect 27834 389494 28454 424938
rect 27834 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 28454 389494
rect 27834 389174 28454 389258
rect 27834 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 28454 389174
rect 27834 353494 28454 388938
rect 27834 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 28454 353494
rect 27834 353174 28454 353258
rect 27834 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 28454 353174
rect 27834 317494 28454 352938
rect 27834 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 28454 317494
rect 27834 317174 28454 317258
rect 27834 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 28454 317174
rect 27834 281494 28454 316938
rect 27834 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 28454 281494
rect 27834 281174 28454 281258
rect 27834 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 28454 281174
rect 27834 245494 28454 280938
rect 27834 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 28454 245494
rect 27834 245174 28454 245258
rect 27834 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 28454 245174
rect 27834 209494 28454 244938
rect 27834 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 28454 209494
rect 27834 209174 28454 209258
rect 27834 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 28454 209174
rect 27834 173494 28454 208938
rect 27834 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 28454 173494
rect 27834 173174 28454 173258
rect 27834 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 28454 173174
rect 27834 137494 28454 172938
rect 27834 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 28454 137494
rect 27834 137174 28454 137258
rect 27834 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 28454 137174
rect 27834 101494 28454 136938
rect 27834 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 28454 101494
rect 27834 101174 28454 101258
rect 27834 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 28454 101174
rect 27834 65494 28454 100938
rect 27834 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 28454 65494
rect 27834 65174 28454 65258
rect 27834 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 28454 65174
rect 27834 29494 28454 64938
rect 27834 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 28454 29494
rect 27834 29174 28454 29258
rect 27834 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 28454 29174
rect 27834 -7066 28454 28938
rect 27834 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 28454 -7066
rect 27834 -7386 28454 -7302
rect 27834 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 28454 -7386
rect 27834 -7654 28454 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 41514 705798 42134 711590
rect 41514 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 42134 705798
rect 41514 705478 42134 705562
rect 41514 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 42134 705478
rect 41514 691174 42134 705242
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -1306 42134 6618
rect 41514 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 42134 -1306
rect 41514 -1626 42134 -1542
rect 41514 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 42134 -1626
rect 41514 -7654 42134 -1862
rect 45234 706758 45854 711590
rect 45234 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 45854 706758
rect 45234 706438 45854 706522
rect 45234 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 45854 706438
rect 45234 694894 45854 706202
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -2266 45854 10338
rect 45234 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 45854 -2266
rect 45234 -2586 45854 -2502
rect 45234 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 45854 -2586
rect 45234 -7654 45854 -2822
rect 48954 707718 49574 711590
rect 48954 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 49574 707718
rect 48954 707398 49574 707482
rect 48954 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 49574 707398
rect 48954 698614 49574 707162
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 48954 -3226 49574 14058
rect 48954 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 49574 -3226
rect 48954 -3546 49574 -3462
rect 48954 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 49574 -3546
rect 48954 -7654 49574 -3782
rect 52674 708678 53294 711590
rect 52674 708442 52706 708678
rect 52942 708442 53026 708678
rect 53262 708442 53294 708678
rect 52674 708358 53294 708442
rect 52674 708122 52706 708358
rect 52942 708122 53026 708358
rect 53262 708122 53294 708358
rect 52674 666334 53294 708122
rect 52674 666098 52706 666334
rect 52942 666098 53026 666334
rect 53262 666098 53294 666334
rect 52674 666014 53294 666098
rect 52674 665778 52706 666014
rect 52942 665778 53026 666014
rect 53262 665778 53294 666014
rect 52674 630334 53294 665778
rect 52674 630098 52706 630334
rect 52942 630098 53026 630334
rect 53262 630098 53294 630334
rect 52674 630014 53294 630098
rect 52674 629778 52706 630014
rect 52942 629778 53026 630014
rect 53262 629778 53294 630014
rect 52674 594334 53294 629778
rect 52674 594098 52706 594334
rect 52942 594098 53026 594334
rect 53262 594098 53294 594334
rect 52674 594014 53294 594098
rect 52674 593778 52706 594014
rect 52942 593778 53026 594014
rect 53262 593778 53294 594014
rect 52674 558334 53294 593778
rect 52674 558098 52706 558334
rect 52942 558098 53026 558334
rect 53262 558098 53294 558334
rect 52674 558014 53294 558098
rect 52674 557778 52706 558014
rect 52942 557778 53026 558014
rect 53262 557778 53294 558014
rect 52674 522334 53294 557778
rect 52674 522098 52706 522334
rect 52942 522098 53026 522334
rect 53262 522098 53294 522334
rect 52674 522014 53294 522098
rect 52674 521778 52706 522014
rect 52942 521778 53026 522014
rect 53262 521778 53294 522014
rect 52674 486334 53294 521778
rect 52674 486098 52706 486334
rect 52942 486098 53026 486334
rect 53262 486098 53294 486334
rect 52674 486014 53294 486098
rect 52674 485778 52706 486014
rect 52942 485778 53026 486014
rect 53262 485778 53294 486014
rect 52674 450334 53294 485778
rect 52674 450098 52706 450334
rect 52942 450098 53026 450334
rect 53262 450098 53294 450334
rect 52674 450014 53294 450098
rect 52674 449778 52706 450014
rect 52942 449778 53026 450014
rect 53262 449778 53294 450014
rect 52674 414334 53294 449778
rect 52674 414098 52706 414334
rect 52942 414098 53026 414334
rect 53262 414098 53294 414334
rect 52674 414014 53294 414098
rect 52674 413778 52706 414014
rect 52942 413778 53026 414014
rect 53262 413778 53294 414014
rect 52674 378334 53294 413778
rect 52674 378098 52706 378334
rect 52942 378098 53026 378334
rect 53262 378098 53294 378334
rect 52674 378014 53294 378098
rect 52674 377778 52706 378014
rect 52942 377778 53026 378014
rect 53262 377778 53294 378014
rect 52674 342334 53294 377778
rect 52674 342098 52706 342334
rect 52942 342098 53026 342334
rect 53262 342098 53294 342334
rect 52674 342014 53294 342098
rect 52674 341778 52706 342014
rect 52942 341778 53026 342014
rect 53262 341778 53294 342014
rect 52674 306334 53294 341778
rect 52674 306098 52706 306334
rect 52942 306098 53026 306334
rect 53262 306098 53294 306334
rect 52674 306014 53294 306098
rect 52674 305778 52706 306014
rect 52942 305778 53026 306014
rect 53262 305778 53294 306014
rect 52674 270334 53294 305778
rect 52674 270098 52706 270334
rect 52942 270098 53026 270334
rect 53262 270098 53294 270334
rect 52674 270014 53294 270098
rect 52674 269778 52706 270014
rect 52942 269778 53026 270014
rect 53262 269778 53294 270014
rect 52674 234334 53294 269778
rect 52674 234098 52706 234334
rect 52942 234098 53026 234334
rect 53262 234098 53294 234334
rect 52674 234014 53294 234098
rect 52674 233778 52706 234014
rect 52942 233778 53026 234014
rect 53262 233778 53294 234014
rect 52674 198334 53294 233778
rect 52674 198098 52706 198334
rect 52942 198098 53026 198334
rect 53262 198098 53294 198334
rect 52674 198014 53294 198098
rect 52674 197778 52706 198014
rect 52942 197778 53026 198014
rect 53262 197778 53294 198014
rect 52674 162334 53294 197778
rect 52674 162098 52706 162334
rect 52942 162098 53026 162334
rect 53262 162098 53294 162334
rect 52674 162014 53294 162098
rect 52674 161778 52706 162014
rect 52942 161778 53026 162014
rect 53262 161778 53294 162014
rect 52674 126334 53294 161778
rect 52674 126098 52706 126334
rect 52942 126098 53026 126334
rect 53262 126098 53294 126334
rect 52674 126014 53294 126098
rect 52674 125778 52706 126014
rect 52942 125778 53026 126014
rect 53262 125778 53294 126014
rect 52674 90334 53294 125778
rect 52674 90098 52706 90334
rect 52942 90098 53026 90334
rect 53262 90098 53294 90334
rect 52674 90014 53294 90098
rect 52674 89778 52706 90014
rect 52942 89778 53026 90014
rect 53262 89778 53294 90014
rect 52674 54334 53294 89778
rect 52674 54098 52706 54334
rect 52942 54098 53026 54334
rect 53262 54098 53294 54334
rect 52674 54014 53294 54098
rect 52674 53778 52706 54014
rect 52942 53778 53026 54014
rect 53262 53778 53294 54014
rect 52674 18334 53294 53778
rect 52674 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 53294 18334
rect 52674 18014 53294 18098
rect 52674 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 53294 18014
rect 52674 -4186 53294 17778
rect 52674 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 53294 -4186
rect 52674 -4506 53294 -4422
rect 52674 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 53294 -4506
rect 52674 -7654 53294 -4742
rect 56394 709638 57014 711590
rect 56394 709402 56426 709638
rect 56662 709402 56746 709638
rect 56982 709402 57014 709638
rect 56394 709318 57014 709402
rect 56394 709082 56426 709318
rect 56662 709082 56746 709318
rect 56982 709082 57014 709318
rect 56394 670054 57014 709082
rect 56394 669818 56426 670054
rect 56662 669818 56746 670054
rect 56982 669818 57014 670054
rect 56394 669734 57014 669818
rect 56394 669498 56426 669734
rect 56662 669498 56746 669734
rect 56982 669498 57014 669734
rect 56394 634054 57014 669498
rect 56394 633818 56426 634054
rect 56662 633818 56746 634054
rect 56982 633818 57014 634054
rect 56394 633734 57014 633818
rect 56394 633498 56426 633734
rect 56662 633498 56746 633734
rect 56982 633498 57014 633734
rect 56394 598054 57014 633498
rect 56394 597818 56426 598054
rect 56662 597818 56746 598054
rect 56982 597818 57014 598054
rect 56394 597734 57014 597818
rect 56394 597498 56426 597734
rect 56662 597498 56746 597734
rect 56982 597498 57014 597734
rect 56394 562054 57014 597498
rect 56394 561818 56426 562054
rect 56662 561818 56746 562054
rect 56982 561818 57014 562054
rect 56394 561734 57014 561818
rect 56394 561498 56426 561734
rect 56662 561498 56746 561734
rect 56982 561498 57014 561734
rect 56394 526054 57014 561498
rect 56394 525818 56426 526054
rect 56662 525818 56746 526054
rect 56982 525818 57014 526054
rect 56394 525734 57014 525818
rect 56394 525498 56426 525734
rect 56662 525498 56746 525734
rect 56982 525498 57014 525734
rect 56394 490054 57014 525498
rect 56394 489818 56426 490054
rect 56662 489818 56746 490054
rect 56982 489818 57014 490054
rect 56394 489734 57014 489818
rect 56394 489498 56426 489734
rect 56662 489498 56746 489734
rect 56982 489498 57014 489734
rect 56394 454054 57014 489498
rect 56394 453818 56426 454054
rect 56662 453818 56746 454054
rect 56982 453818 57014 454054
rect 56394 453734 57014 453818
rect 56394 453498 56426 453734
rect 56662 453498 56746 453734
rect 56982 453498 57014 453734
rect 56394 418054 57014 453498
rect 56394 417818 56426 418054
rect 56662 417818 56746 418054
rect 56982 417818 57014 418054
rect 56394 417734 57014 417818
rect 56394 417498 56426 417734
rect 56662 417498 56746 417734
rect 56982 417498 57014 417734
rect 56394 382054 57014 417498
rect 56394 381818 56426 382054
rect 56662 381818 56746 382054
rect 56982 381818 57014 382054
rect 56394 381734 57014 381818
rect 56394 381498 56426 381734
rect 56662 381498 56746 381734
rect 56982 381498 57014 381734
rect 56394 346054 57014 381498
rect 56394 345818 56426 346054
rect 56662 345818 56746 346054
rect 56982 345818 57014 346054
rect 56394 345734 57014 345818
rect 56394 345498 56426 345734
rect 56662 345498 56746 345734
rect 56982 345498 57014 345734
rect 56394 310054 57014 345498
rect 56394 309818 56426 310054
rect 56662 309818 56746 310054
rect 56982 309818 57014 310054
rect 56394 309734 57014 309818
rect 56394 309498 56426 309734
rect 56662 309498 56746 309734
rect 56982 309498 57014 309734
rect 56394 274054 57014 309498
rect 56394 273818 56426 274054
rect 56662 273818 56746 274054
rect 56982 273818 57014 274054
rect 56394 273734 57014 273818
rect 56394 273498 56426 273734
rect 56662 273498 56746 273734
rect 56982 273498 57014 273734
rect 56394 238054 57014 273498
rect 56394 237818 56426 238054
rect 56662 237818 56746 238054
rect 56982 237818 57014 238054
rect 56394 237734 57014 237818
rect 56394 237498 56426 237734
rect 56662 237498 56746 237734
rect 56982 237498 57014 237734
rect 56394 202054 57014 237498
rect 56394 201818 56426 202054
rect 56662 201818 56746 202054
rect 56982 201818 57014 202054
rect 56394 201734 57014 201818
rect 56394 201498 56426 201734
rect 56662 201498 56746 201734
rect 56982 201498 57014 201734
rect 56394 166054 57014 201498
rect 56394 165818 56426 166054
rect 56662 165818 56746 166054
rect 56982 165818 57014 166054
rect 56394 165734 57014 165818
rect 56394 165498 56426 165734
rect 56662 165498 56746 165734
rect 56982 165498 57014 165734
rect 56394 130054 57014 165498
rect 56394 129818 56426 130054
rect 56662 129818 56746 130054
rect 56982 129818 57014 130054
rect 56394 129734 57014 129818
rect 56394 129498 56426 129734
rect 56662 129498 56746 129734
rect 56982 129498 57014 129734
rect 56394 94054 57014 129498
rect 56394 93818 56426 94054
rect 56662 93818 56746 94054
rect 56982 93818 57014 94054
rect 56394 93734 57014 93818
rect 56394 93498 56426 93734
rect 56662 93498 56746 93734
rect 56982 93498 57014 93734
rect 56394 58054 57014 93498
rect 56394 57818 56426 58054
rect 56662 57818 56746 58054
rect 56982 57818 57014 58054
rect 56394 57734 57014 57818
rect 56394 57498 56426 57734
rect 56662 57498 56746 57734
rect 56982 57498 57014 57734
rect 56394 22054 57014 57498
rect 56394 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 57014 22054
rect 56394 21734 57014 21818
rect 56394 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 57014 21734
rect 56394 -5146 57014 21498
rect 56394 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 57014 -5146
rect 56394 -5466 57014 -5382
rect 56394 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 57014 -5466
rect 56394 -7654 57014 -5702
rect 60114 710598 60734 711590
rect 60114 710362 60146 710598
rect 60382 710362 60466 710598
rect 60702 710362 60734 710598
rect 60114 710278 60734 710362
rect 60114 710042 60146 710278
rect 60382 710042 60466 710278
rect 60702 710042 60734 710278
rect 60114 673774 60734 710042
rect 60114 673538 60146 673774
rect 60382 673538 60466 673774
rect 60702 673538 60734 673774
rect 60114 673454 60734 673538
rect 60114 673218 60146 673454
rect 60382 673218 60466 673454
rect 60702 673218 60734 673454
rect 60114 637774 60734 673218
rect 60114 637538 60146 637774
rect 60382 637538 60466 637774
rect 60702 637538 60734 637774
rect 60114 637454 60734 637538
rect 60114 637218 60146 637454
rect 60382 637218 60466 637454
rect 60702 637218 60734 637454
rect 60114 601774 60734 637218
rect 60114 601538 60146 601774
rect 60382 601538 60466 601774
rect 60702 601538 60734 601774
rect 60114 601454 60734 601538
rect 60114 601218 60146 601454
rect 60382 601218 60466 601454
rect 60702 601218 60734 601454
rect 60114 565774 60734 601218
rect 60114 565538 60146 565774
rect 60382 565538 60466 565774
rect 60702 565538 60734 565774
rect 60114 565454 60734 565538
rect 60114 565218 60146 565454
rect 60382 565218 60466 565454
rect 60702 565218 60734 565454
rect 60114 529774 60734 565218
rect 60114 529538 60146 529774
rect 60382 529538 60466 529774
rect 60702 529538 60734 529774
rect 60114 529454 60734 529538
rect 60114 529218 60146 529454
rect 60382 529218 60466 529454
rect 60702 529218 60734 529454
rect 60114 493774 60734 529218
rect 60114 493538 60146 493774
rect 60382 493538 60466 493774
rect 60702 493538 60734 493774
rect 60114 493454 60734 493538
rect 60114 493218 60146 493454
rect 60382 493218 60466 493454
rect 60702 493218 60734 493454
rect 60114 457774 60734 493218
rect 60114 457538 60146 457774
rect 60382 457538 60466 457774
rect 60702 457538 60734 457774
rect 60114 457454 60734 457538
rect 60114 457218 60146 457454
rect 60382 457218 60466 457454
rect 60702 457218 60734 457454
rect 60114 421774 60734 457218
rect 60114 421538 60146 421774
rect 60382 421538 60466 421774
rect 60702 421538 60734 421774
rect 60114 421454 60734 421538
rect 60114 421218 60146 421454
rect 60382 421218 60466 421454
rect 60702 421218 60734 421454
rect 60114 385774 60734 421218
rect 60114 385538 60146 385774
rect 60382 385538 60466 385774
rect 60702 385538 60734 385774
rect 60114 385454 60734 385538
rect 60114 385218 60146 385454
rect 60382 385218 60466 385454
rect 60702 385218 60734 385454
rect 60114 349774 60734 385218
rect 60114 349538 60146 349774
rect 60382 349538 60466 349774
rect 60702 349538 60734 349774
rect 60114 349454 60734 349538
rect 60114 349218 60146 349454
rect 60382 349218 60466 349454
rect 60702 349218 60734 349454
rect 60114 313774 60734 349218
rect 60114 313538 60146 313774
rect 60382 313538 60466 313774
rect 60702 313538 60734 313774
rect 60114 313454 60734 313538
rect 60114 313218 60146 313454
rect 60382 313218 60466 313454
rect 60702 313218 60734 313454
rect 60114 277774 60734 313218
rect 60114 277538 60146 277774
rect 60382 277538 60466 277774
rect 60702 277538 60734 277774
rect 60114 277454 60734 277538
rect 60114 277218 60146 277454
rect 60382 277218 60466 277454
rect 60702 277218 60734 277454
rect 60114 241774 60734 277218
rect 60114 241538 60146 241774
rect 60382 241538 60466 241774
rect 60702 241538 60734 241774
rect 60114 241454 60734 241538
rect 60114 241218 60146 241454
rect 60382 241218 60466 241454
rect 60702 241218 60734 241454
rect 60114 205774 60734 241218
rect 60114 205538 60146 205774
rect 60382 205538 60466 205774
rect 60702 205538 60734 205774
rect 60114 205454 60734 205538
rect 60114 205218 60146 205454
rect 60382 205218 60466 205454
rect 60702 205218 60734 205454
rect 60114 169774 60734 205218
rect 60114 169538 60146 169774
rect 60382 169538 60466 169774
rect 60702 169538 60734 169774
rect 60114 169454 60734 169538
rect 60114 169218 60146 169454
rect 60382 169218 60466 169454
rect 60702 169218 60734 169454
rect 60114 133774 60734 169218
rect 60114 133538 60146 133774
rect 60382 133538 60466 133774
rect 60702 133538 60734 133774
rect 60114 133454 60734 133538
rect 60114 133218 60146 133454
rect 60382 133218 60466 133454
rect 60702 133218 60734 133454
rect 60114 97774 60734 133218
rect 60114 97538 60146 97774
rect 60382 97538 60466 97774
rect 60702 97538 60734 97774
rect 60114 97454 60734 97538
rect 60114 97218 60146 97454
rect 60382 97218 60466 97454
rect 60702 97218 60734 97454
rect 60114 61774 60734 97218
rect 60114 61538 60146 61774
rect 60382 61538 60466 61774
rect 60702 61538 60734 61774
rect 60114 61454 60734 61538
rect 60114 61218 60146 61454
rect 60382 61218 60466 61454
rect 60702 61218 60734 61454
rect 60114 25774 60734 61218
rect 60114 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 60734 25774
rect 60114 25454 60734 25538
rect 60114 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 60734 25454
rect 60114 -6106 60734 25218
rect 60114 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 60734 -6106
rect 60114 -6426 60734 -6342
rect 60114 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 60734 -6426
rect 60114 -7654 60734 -6662
rect 63834 711558 64454 711590
rect 63834 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 64454 711558
rect 63834 711238 64454 711322
rect 63834 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 64454 711238
rect 63834 677494 64454 711002
rect 63834 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 64454 677494
rect 63834 677174 64454 677258
rect 63834 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 64454 677174
rect 63834 641494 64454 676938
rect 63834 641258 63866 641494
rect 64102 641258 64186 641494
rect 64422 641258 64454 641494
rect 63834 641174 64454 641258
rect 63834 640938 63866 641174
rect 64102 640938 64186 641174
rect 64422 640938 64454 641174
rect 63834 605494 64454 640938
rect 63834 605258 63866 605494
rect 64102 605258 64186 605494
rect 64422 605258 64454 605494
rect 63834 605174 64454 605258
rect 63834 604938 63866 605174
rect 64102 604938 64186 605174
rect 64422 604938 64454 605174
rect 63834 569494 64454 604938
rect 63834 569258 63866 569494
rect 64102 569258 64186 569494
rect 64422 569258 64454 569494
rect 63834 569174 64454 569258
rect 63834 568938 63866 569174
rect 64102 568938 64186 569174
rect 64422 568938 64454 569174
rect 63834 533494 64454 568938
rect 63834 533258 63866 533494
rect 64102 533258 64186 533494
rect 64422 533258 64454 533494
rect 63834 533174 64454 533258
rect 63834 532938 63866 533174
rect 64102 532938 64186 533174
rect 64422 532938 64454 533174
rect 63834 497494 64454 532938
rect 63834 497258 63866 497494
rect 64102 497258 64186 497494
rect 64422 497258 64454 497494
rect 63834 497174 64454 497258
rect 63834 496938 63866 497174
rect 64102 496938 64186 497174
rect 64422 496938 64454 497174
rect 63834 461494 64454 496938
rect 63834 461258 63866 461494
rect 64102 461258 64186 461494
rect 64422 461258 64454 461494
rect 63834 461174 64454 461258
rect 63834 460938 63866 461174
rect 64102 460938 64186 461174
rect 64422 460938 64454 461174
rect 63834 425494 64454 460938
rect 63834 425258 63866 425494
rect 64102 425258 64186 425494
rect 64422 425258 64454 425494
rect 63834 425174 64454 425258
rect 63834 424938 63866 425174
rect 64102 424938 64186 425174
rect 64422 424938 64454 425174
rect 63834 389494 64454 424938
rect 63834 389258 63866 389494
rect 64102 389258 64186 389494
rect 64422 389258 64454 389494
rect 63834 389174 64454 389258
rect 63834 388938 63866 389174
rect 64102 388938 64186 389174
rect 64422 388938 64454 389174
rect 63834 353494 64454 388938
rect 63834 353258 63866 353494
rect 64102 353258 64186 353494
rect 64422 353258 64454 353494
rect 63834 353174 64454 353258
rect 63834 352938 63866 353174
rect 64102 352938 64186 353174
rect 64422 352938 64454 353174
rect 63834 317494 64454 352938
rect 63834 317258 63866 317494
rect 64102 317258 64186 317494
rect 64422 317258 64454 317494
rect 63834 317174 64454 317258
rect 63834 316938 63866 317174
rect 64102 316938 64186 317174
rect 64422 316938 64454 317174
rect 63834 281494 64454 316938
rect 63834 281258 63866 281494
rect 64102 281258 64186 281494
rect 64422 281258 64454 281494
rect 63834 281174 64454 281258
rect 63834 280938 63866 281174
rect 64102 280938 64186 281174
rect 64422 280938 64454 281174
rect 63834 245494 64454 280938
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 68323 252924 68389 252925
rect 68323 252860 68324 252924
rect 68388 252860 68389 252924
rect 68323 252859 68389 252860
rect 63834 245258 63866 245494
rect 64102 245258 64186 245494
rect 64422 245258 64454 245494
rect 63834 245174 64454 245258
rect 63834 244938 63866 245174
rect 64102 244938 64186 245174
rect 64422 244938 64454 245174
rect 63834 209494 64454 244938
rect 67219 241636 67285 241637
rect 67219 241572 67220 241636
rect 67284 241572 67285 241636
rect 67219 241571 67285 241572
rect 63834 209258 63866 209494
rect 64102 209258 64186 209494
rect 64422 209258 64454 209494
rect 63834 209174 64454 209258
rect 63834 208938 63866 209174
rect 64102 208938 64186 209174
rect 64422 208938 64454 209174
rect 63834 173494 64454 208938
rect 63834 173258 63866 173494
rect 64102 173258 64186 173494
rect 64422 173258 64454 173494
rect 63834 173174 64454 173258
rect 63834 172938 63866 173174
rect 64102 172938 64186 173174
rect 64422 172938 64454 173174
rect 63834 137494 64454 172938
rect 63834 137258 63866 137494
rect 64102 137258 64186 137494
rect 64422 137258 64454 137494
rect 63834 137174 64454 137258
rect 63834 136938 63866 137174
rect 64102 136938 64186 137174
rect 64422 136938 64454 137174
rect 63834 101494 64454 136938
rect 67222 112437 67282 241571
rect 68326 239597 68386 252859
rect 68691 252788 68757 252789
rect 68691 252724 68692 252788
rect 68756 252724 68757 252788
rect 68691 252723 68757 252724
rect 68507 252652 68573 252653
rect 68507 252588 68508 252652
rect 68572 252588 68573 252652
rect 68507 252587 68573 252588
rect 68323 239596 68389 239597
rect 68323 239532 68324 239596
rect 68388 239532 68389 239596
rect 68323 239531 68389 239532
rect 68510 238917 68570 252587
rect 68507 238916 68573 238917
rect 68507 238852 68508 238916
rect 68572 238852 68573 238916
rect 68507 238851 68573 238852
rect 68694 232661 68754 252723
rect 69059 251836 69125 251837
rect 69059 251772 69060 251836
rect 69124 251772 69125 251836
rect 69059 251771 69125 251772
rect 68875 248300 68941 248301
rect 68875 248236 68876 248300
rect 68940 248236 68941 248300
rect 68875 248235 68941 248236
rect 68691 232660 68757 232661
rect 68691 232596 68692 232660
rect 68756 232596 68757 232660
rect 68691 232595 68757 232596
rect 68691 210220 68757 210221
rect 68691 210156 68692 210220
rect 68756 210156 68757 210220
rect 68691 210155 68757 210156
rect 68507 205596 68573 205597
rect 68507 205532 68508 205596
rect 68572 205532 68573 205596
rect 68507 205531 68573 205532
rect 68323 203420 68389 203421
rect 68323 203356 68324 203420
rect 68388 203356 68389 203420
rect 68323 203355 68389 203356
rect 67403 200156 67469 200157
rect 67403 200092 67404 200156
rect 67468 200092 67469 200156
rect 67403 200091 67469 200092
rect 67219 112436 67285 112437
rect 67219 112372 67220 112436
rect 67284 112372 67285 112436
rect 67219 112371 67285 112372
rect 67222 102101 67282 112371
rect 67219 102100 67285 102101
rect 67219 102036 67220 102100
rect 67284 102036 67285 102100
rect 67219 102035 67285 102036
rect 63834 101258 63866 101494
rect 64102 101258 64186 101494
rect 64422 101258 64454 101494
rect 63834 101174 64454 101258
rect 63834 100938 63866 101174
rect 64102 100938 64186 101174
rect 64422 100938 64454 101174
rect 63834 65494 64454 100938
rect 67406 75717 67466 200091
rect 68326 174045 68386 203355
rect 68510 177309 68570 205531
rect 68694 198797 68754 210155
rect 68691 198796 68757 198797
rect 68691 198732 68692 198796
rect 68756 198732 68757 198796
rect 68691 198731 68757 198732
rect 68507 177308 68573 177309
rect 68507 177244 68508 177308
rect 68572 177244 68573 177308
rect 68507 177243 68573 177244
rect 68323 174044 68389 174045
rect 68323 173980 68324 174044
rect 68388 173980 68389 174044
rect 68323 173979 68389 173980
rect 67403 75716 67469 75717
rect 67403 75652 67404 75716
rect 67468 75652 67469 75716
rect 67403 75651 67469 75652
rect 68326 73269 68386 173979
rect 68510 74085 68570 177243
rect 68878 117333 68938 248235
rect 68875 117332 68941 117333
rect 68875 117268 68876 117332
rect 68940 117268 68941 117332
rect 68875 117267 68941 117268
rect 69062 110941 69122 251771
rect 73794 249436 74414 254898
rect 77514 705798 78134 711590
rect 77514 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 78134 705798
rect 77514 705478 78134 705562
rect 77514 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 78134 705478
rect 77514 691174 78134 705242
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 74208 219454 74528 219486
rect 74208 219218 74250 219454
rect 74486 219218 74528 219454
rect 74208 219134 74528 219218
rect 74208 218898 74250 219134
rect 74486 218898 74528 219134
rect 74208 218866 74528 218898
rect 70715 209540 70781 209541
rect 70715 209476 70716 209540
rect 70780 209476 70781 209540
rect 70715 209475 70781 209476
rect 69243 207500 69309 207501
rect 69243 207436 69244 207500
rect 69308 207436 69309 207500
rect 69243 207435 69309 207436
rect 69246 200157 69306 207435
rect 70718 205650 70778 209475
rect 70534 205590 70778 205650
rect 69795 204916 69861 204917
rect 69795 204852 69796 204916
rect 69860 204852 69861 204916
rect 69795 204851 69861 204852
rect 69611 201244 69677 201245
rect 69611 201180 69612 201244
rect 69676 201180 69677 201244
rect 69611 201179 69677 201180
rect 69243 200156 69309 200157
rect 69243 200092 69244 200156
rect 69308 200092 69309 200156
rect 69243 200091 69309 200092
rect 69246 179349 69306 200091
rect 69614 189005 69674 201179
rect 69798 194581 69858 204851
rect 70163 200292 70229 200293
rect 70163 200228 70164 200292
rect 70228 200290 70229 200292
rect 70534 200290 70594 205590
rect 70228 200230 70594 200290
rect 70228 200228 70229 200230
rect 70163 200227 70229 200228
rect 70534 195990 70594 200230
rect 70534 195930 71146 195990
rect 69795 194580 69861 194581
rect 69795 194516 69796 194580
rect 69860 194516 69861 194580
rect 69795 194515 69861 194516
rect 69611 189004 69677 189005
rect 69611 188940 69612 189004
rect 69676 188940 69677 189004
rect 69611 188939 69677 188940
rect 71086 180845 71146 195930
rect 73794 183454 74414 200068
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 71267 180980 71333 180981
rect 71267 180916 71268 180980
rect 71332 180916 71333 180980
rect 71267 180915 71333 180916
rect 71083 180844 71149 180845
rect 71083 180780 71084 180844
rect 71148 180780 71149 180844
rect 71083 180779 71149 180780
rect 69243 179348 69309 179349
rect 69243 179284 69244 179348
rect 69308 179284 69309 179348
rect 69243 179283 69309 179284
rect 71270 178125 71330 180915
rect 71267 178124 71333 178125
rect 71267 178060 71268 178124
rect 71332 178060 71333 178124
rect 71267 178059 71333 178060
rect 69243 175948 69309 175949
rect 69243 175884 69244 175948
rect 69308 175884 69309 175948
rect 69243 175883 69309 175884
rect 69059 110940 69125 110941
rect 69059 110876 69060 110940
rect 69124 110876 69125 110940
rect 69059 110875 69125 110876
rect 69059 84964 69125 84965
rect 69059 84900 69060 84964
rect 69124 84900 69125 84964
rect 69059 84899 69125 84900
rect 68691 83604 68757 83605
rect 68691 83540 68692 83604
rect 68756 83540 68757 83604
rect 68691 83539 68757 83540
rect 68507 74084 68573 74085
rect 68507 74020 68508 74084
rect 68572 74020 68573 74084
rect 68507 74019 68573 74020
rect 68323 73268 68389 73269
rect 68323 73204 68324 73268
rect 68388 73204 68389 73268
rect 68323 73203 68389 73204
rect 68694 69597 68754 83539
rect 68875 75716 68941 75717
rect 68875 75652 68876 75716
rect 68940 75652 68941 75716
rect 68875 75651 68941 75652
rect 68691 69596 68757 69597
rect 68691 69532 68692 69596
rect 68756 69532 68757 69596
rect 68691 69531 68757 69532
rect 68878 69461 68938 75651
rect 69062 69869 69122 84899
rect 69246 73405 69306 175883
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 70531 112572 70597 112573
rect 70531 112508 70532 112572
rect 70596 112508 70597 112572
rect 70531 112507 70597 112508
rect 69427 112028 69493 112029
rect 69427 111964 69428 112028
rect 69492 111964 69493 112028
rect 69427 111963 69493 111964
rect 69430 92581 69490 111963
rect 70163 111892 70229 111893
rect 70163 111828 70164 111892
rect 70228 111828 70229 111892
rect 70163 111827 70229 111828
rect 70166 111349 70226 111827
rect 70163 111348 70229 111349
rect 70163 111284 70164 111348
rect 70228 111284 70229 111348
rect 70163 111283 70229 111284
rect 70534 109050 70594 112507
rect 70350 108990 70594 109050
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 70350 108901 70410 108990
rect 70347 108900 70413 108901
rect 70347 108836 70348 108900
rect 70412 108836 70413 108900
rect 70347 108835 70413 108836
rect 69427 92580 69493 92581
rect 69427 92516 69428 92580
rect 69492 92516 69493 92580
rect 69427 92515 69493 92516
rect 73794 75454 74414 110898
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 81234 706758 81854 711590
rect 81234 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 81854 706758
rect 81234 706438 81854 706522
rect 81234 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 81854 706438
rect 81234 694894 81854 706202
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 118894 81854 154338
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 69243 73404 69309 73405
rect 69243 73340 69244 73404
rect 69308 73340 69309 73404
rect 69243 73339 69309 73340
rect 70531 73268 70597 73269
rect 70531 73204 70532 73268
rect 70596 73204 70597 73268
rect 70531 73203 70597 73204
rect 70534 70005 70594 73203
rect 70531 70004 70597 70005
rect 70531 69940 70532 70004
rect 70596 69940 70597 70004
rect 70531 69939 70597 69940
rect 69059 69868 69125 69869
rect 69059 69804 69060 69868
rect 69124 69804 69125 69868
rect 69059 69803 69125 69804
rect 68875 69460 68941 69461
rect 68875 69396 68876 69460
rect 68940 69396 68941 69460
rect 68875 69395 68941 69396
rect 63834 65258 63866 65494
rect 64102 65258 64186 65494
rect 64422 65258 64454 65494
rect 63834 65174 64454 65258
rect 63834 64938 63866 65174
rect 64102 64938 64186 65174
rect 64422 64938 64454 65174
rect 63834 29494 64454 64938
rect 63834 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 64454 29494
rect 63834 29174 64454 29258
rect 63834 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 64454 29174
rect 63834 -7066 64454 28938
rect 63834 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 64454 -7066
rect 63834 -7386 64454 -7302
rect 63834 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 64454 -7386
rect 63834 -7654 64454 -7622
rect 73794 39454 74414 74898
rect 75164 75454 75484 75486
rect 75164 75218 75206 75454
rect 75442 75218 75484 75454
rect 75164 75134 75484 75218
rect 75164 74898 75206 75134
rect 75442 74898 75484 75134
rect 75164 74866 75484 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 77514 43174 78134 78618
rect 79384 79174 79704 79206
rect 79384 78938 79426 79174
rect 79662 78938 79704 79174
rect 79384 78854 79704 78938
rect 79384 78618 79426 78854
rect 79662 78618 79704 78854
rect 79384 78586 79704 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -1306 78134 6618
rect 77514 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 78134 -1306
rect 77514 -1626 78134 -1542
rect 77514 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 78134 -1626
rect 77514 -7654 78134 -1862
rect 81234 46894 81854 82338
rect 84954 707718 85574 711590
rect 84954 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 85574 707718
rect 84954 707398 85574 707482
rect 84954 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 85574 707398
rect 84954 698614 85574 707162
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 88674 708678 89294 711590
rect 88674 708442 88706 708678
rect 88942 708442 89026 708678
rect 89262 708442 89294 708678
rect 88674 708358 89294 708442
rect 88674 708122 88706 708358
rect 88942 708122 89026 708358
rect 89262 708122 89294 708358
rect 88674 666334 89294 708122
rect 88674 666098 88706 666334
rect 88942 666098 89026 666334
rect 89262 666098 89294 666334
rect 88674 666014 89294 666098
rect 88674 665778 88706 666014
rect 88942 665778 89026 666014
rect 89262 665778 89294 666014
rect 88674 630334 89294 665778
rect 88674 630098 88706 630334
rect 88942 630098 89026 630334
rect 89262 630098 89294 630334
rect 88674 630014 89294 630098
rect 88674 629778 88706 630014
rect 88942 629778 89026 630014
rect 89262 629778 89294 630014
rect 88674 594334 89294 629778
rect 88674 594098 88706 594334
rect 88942 594098 89026 594334
rect 89262 594098 89294 594334
rect 88674 594014 89294 594098
rect 88674 593778 88706 594014
rect 88942 593778 89026 594014
rect 89262 593778 89294 594014
rect 88674 558334 89294 593778
rect 88674 558098 88706 558334
rect 88942 558098 89026 558334
rect 89262 558098 89294 558334
rect 88674 558014 89294 558098
rect 88674 557778 88706 558014
rect 88942 557778 89026 558014
rect 89262 557778 89294 558014
rect 88674 522334 89294 557778
rect 88674 522098 88706 522334
rect 88942 522098 89026 522334
rect 89262 522098 89294 522334
rect 88674 522014 89294 522098
rect 88674 521778 88706 522014
rect 88942 521778 89026 522014
rect 89262 521778 89294 522014
rect 88674 486334 89294 521778
rect 88674 486098 88706 486334
rect 88942 486098 89026 486334
rect 89262 486098 89294 486334
rect 88674 486014 89294 486098
rect 88674 485778 88706 486014
rect 88942 485778 89026 486014
rect 89262 485778 89294 486014
rect 88674 450334 89294 485778
rect 88674 450098 88706 450334
rect 88942 450098 89026 450334
rect 89262 450098 89294 450334
rect 88674 450014 89294 450098
rect 88674 449778 88706 450014
rect 88942 449778 89026 450014
rect 89262 449778 89294 450014
rect 88674 414334 89294 449778
rect 88674 414098 88706 414334
rect 88942 414098 89026 414334
rect 89262 414098 89294 414334
rect 88674 414014 89294 414098
rect 88674 413778 88706 414014
rect 88942 413778 89026 414014
rect 89262 413778 89294 414014
rect 88674 378334 89294 413778
rect 88674 378098 88706 378334
rect 88942 378098 89026 378334
rect 89262 378098 89294 378334
rect 88674 378014 89294 378098
rect 88674 377778 88706 378014
rect 88942 377778 89026 378014
rect 89262 377778 89294 378014
rect 88674 342334 89294 377778
rect 88674 342098 88706 342334
rect 88942 342098 89026 342334
rect 89262 342098 89294 342334
rect 88674 342014 89294 342098
rect 88674 341778 88706 342014
rect 88942 341778 89026 342014
rect 89262 341778 89294 342014
rect 88674 306334 89294 341778
rect 88674 306098 88706 306334
rect 88942 306098 89026 306334
rect 89262 306098 89294 306334
rect 88674 306014 89294 306098
rect 88674 305778 88706 306014
rect 88942 305778 89026 306014
rect 89262 305778 89294 306014
rect 88674 270334 89294 305778
rect 88674 270098 88706 270334
rect 88942 270098 89026 270334
rect 89262 270098 89294 270334
rect 88674 270014 89294 270098
rect 88674 269778 88706 270014
rect 88942 269778 89026 270014
rect 89262 269778 89294 270014
rect 88674 249081 89294 269778
rect 92394 709638 93014 711590
rect 92394 709402 92426 709638
rect 92662 709402 92746 709638
rect 92982 709402 93014 709638
rect 92394 709318 93014 709402
rect 92394 709082 92426 709318
rect 92662 709082 92746 709318
rect 92982 709082 93014 709318
rect 92394 670054 93014 709082
rect 92394 669818 92426 670054
rect 92662 669818 92746 670054
rect 92982 669818 93014 670054
rect 92394 669734 93014 669818
rect 92394 669498 92426 669734
rect 92662 669498 92746 669734
rect 92982 669498 93014 669734
rect 92394 634054 93014 669498
rect 92394 633818 92426 634054
rect 92662 633818 92746 634054
rect 92982 633818 93014 634054
rect 92394 633734 93014 633818
rect 92394 633498 92426 633734
rect 92662 633498 92746 633734
rect 92982 633498 93014 633734
rect 92394 598054 93014 633498
rect 92394 597818 92426 598054
rect 92662 597818 92746 598054
rect 92982 597818 93014 598054
rect 92394 597734 93014 597818
rect 92394 597498 92426 597734
rect 92662 597498 92746 597734
rect 92982 597498 93014 597734
rect 92394 562054 93014 597498
rect 92394 561818 92426 562054
rect 92662 561818 92746 562054
rect 92982 561818 93014 562054
rect 92394 561734 93014 561818
rect 92394 561498 92426 561734
rect 92662 561498 92746 561734
rect 92982 561498 93014 561734
rect 92394 526054 93014 561498
rect 92394 525818 92426 526054
rect 92662 525818 92746 526054
rect 92982 525818 93014 526054
rect 92394 525734 93014 525818
rect 92394 525498 92426 525734
rect 92662 525498 92746 525734
rect 92982 525498 93014 525734
rect 92394 490054 93014 525498
rect 92394 489818 92426 490054
rect 92662 489818 92746 490054
rect 92982 489818 93014 490054
rect 92394 489734 93014 489818
rect 92394 489498 92426 489734
rect 92662 489498 92746 489734
rect 92982 489498 93014 489734
rect 92394 454054 93014 489498
rect 92394 453818 92426 454054
rect 92662 453818 92746 454054
rect 92982 453818 93014 454054
rect 92394 453734 93014 453818
rect 92394 453498 92426 453734
rect 92662 453498 92746 453734
rect 92982 453498 93014 453734
rect 92394 418054 93014 453498
rect 92394 417818 92426 418054
rect 92662 417818 92746 418054
rect 92982 417818 93014 418054
rect 92394 417734 93014 417818
rect 92394 417498 92426 417734
rect 92662 417498 92746 417734
rect 92982 417498 93014 417734
rect 92394 382054 93014 417498
rect 92394 381818 92426 382054
rect 92662 381818 92746 382054
rect 92982 381818 93014 382054
rect 92394 381734 93014 381818
rect 92394 381498 92426 381734
rect 92662 381498 92746 381734
rect 92982 381498 93014 381734
rect 92394 346054 93014 381498
rect 92394 345818 92426 346054
rect 92662 345818 92746 346054
rect 92982 345818 93014 346054
rect 92394 345734 93014 345818
rect 92394 345498 92426 345734
rect 92662 345498 92746 345734
rect 92982 345498 93014 345734
rect 92394 310054 93014 345498
rect 92394 309818 92426 310054
rect 92662 309818 92746 310054
rect 92982 309818 93014 310054
rect 92394 309734 93014 309818
rect 92394 309498 92426 309734
rect 92662 309498 92746 309734
rect 92982 309498 93014 309734
rect 92394 274054 93014 309498
rect 92394 273818 92426 274054
rect 92662 273818 92746 274054
rect 92982 273818 93014 274054
rect 92394 273734 93014 273818
rect 92394 273498 92426 273734
rect 92662 273498 92746 273734
rect 92982 273498 93014 273734
rect 92394 249081 93014 273498
rect 96114 710598 96734 711590
rect 96114 710362 96146 710598
rect 96382 710362 96466 710598
rect 96702 710362 96734 710598
rect 96114 710278 96734 710362
rect 96114 710042 96146 710278
rect 96382 710042 96466 710278
rect 96702 710042 96734 710278
rect 96114 673774 96734 710042
rect 96114 673538 96146 673774
rect 96382 673538 96466 673774
rect 96702 673538 96734 673774
rect 96114 673454 96734 673538
rect 96114 673218 96146 673454
rect 96382 673218 96466 673454
rect 96702 673218 96734 673454
rect 96114 637774 96734 673218
rect 96114 637538 96146 637774
rect 96382 637538 96466 637774
rect 96702 637538 96734 637774
rect 96114 637454 96734 637538
rect 96114 637218 96146 637454
rect 96382 637218 96466 637454
rect 96702 637218 96734 637454
rect 96114 601774 96734 637218
rect 96114 601538 96146 601774
rect 96382 601538 96466 601774
rect 96702 601538 96734 601774
rect 96114 601454 96734 601538
rect 96114 601218 96146 601454
rect 96382 601218 96466 601454
rect 96702 601218 96734 601454
rect 96114 565774 96734 601218
rect 96114 565538 96146 565774
rect 96382 565538 96466 565774
rect 96702 565538 96734 565774
rect 96114 565454 96734 565538
rect 96114 565218 96146 565454
rect 96382 565218 96466 565454
rect 96702 565218 96734 565454
rect 96114 529774 96734 565218
rect 96114 529538 96146 529774
rect 96382 529538 96466 529774
rect 96702 529538 96734 529774
rect 96114 529454 96734 529538
rect 96114 529218 96146 529454
rect 96382 529218 96466 529454
rect 96702 529218 96734 529454
rect 96114 493774 96734 529218
rect 96114 493538 96146 493774
rect 96382 493538 96466 493774
rect 96702 493538 96734 493774
rect 96114 493454 96734 493538
rect 96114 493218 96146 493454
rect 96382 493218 96466 493454
rect 96702 493218 96734 493454
rect 96114 457774 96734 493218
rect 96114 457538 96146 457774
rect 96382 457538 96466 457774
rect 96702 457538 96734 457774
rect 96114 457454 96734 457538
rect 96114 457218 96146 457454
rect 96382 457218 96466 457454
rect 96702 457218 96734 457454
rect 96114 421774 96734 457218
rect 96114 421538 96146 421774
rect 96382 421538 96466 421774
rect 96702 421538 96734 421774
rect 96114 421454 96734 421538
rect 96114 421218 96146 421454
rect 96382 421218 96466 421454
rect 96702 421218 96734 421454
rect 96114 385774 96734 421218
rect 96114 385538 96146 385774
rect 96382 385538 96466 385774
rect 96702 385538 96734 385774
rect 96114 385454 96734 385538
rect 96114 385218 96146 385454
rect 96382 385218 96466 385454
rect 96702 385218 96734 385454
rect 96114 349774 96734 385218
rect 96114 349538 96146 349774
rect 96382 349538 96466 349774
rect 96702 349538 96734 349774
rect 96114 349454 96734 349538
rect 96114 349218 96146 349454
rect 96382 349218 96466 349454
rect 96702 349218 96734 349454
rect 96114 313774 96734 349218
rect 96114 313538 96146 313774
rect 96382 313538 96466 313774
rect 96702 313538 96734 313774
rect 96114 313454 96734 313538
rect 96114 313218 96146 313454
rect 96382 313218 96466 313454
rect 96702 313218 96734 313454
rect 96114 277774 96734 313218
rect 96114 277538 96146 277774
rect 96382 277538 96466 277774
rect 96702 277538 96734 277774
rect 96114 277454 96734 277538
rect 96114 277218 96146 277454
rect 96382 277218 96466 277454
rect 96702 277218 96734 277454
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 96114 241774 96734 277218
rect 96114 241538 96146 241774
rect 96382 241538 96466 241774
rect 96702 241538 96734 241774
rect 96114 241454 96734 241538
rect 96114 241218 96146 241454
rect 96382 241218 96466 241454
rect 96702 241218 96734 241454
rect 89568 223174 89888 223206
rect 89568 222938 89610 223174
rect 89846 222938 89888 223174
rect 89568 222854 89888 222938
rect 89568 222618 89610 222854
rect 89846 222618 89888 222854
rect 89568 222586 89888 222618
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 122614 85574 158058
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 83605 75454 83925 75486
rect 83605 75218 83647 75454
rect 83883 75218 83925 75454
rect 83605 75134 83925 75218
rect 83605 74898 83647 75134
rect 83883 74898 83925 75134
rect 83605 74866 83925 74898
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -2266 81854 10338
rect 81234 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 81854 -2266
rect 81234 -2586 81854 -2502
rect 81234 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 81854 -2586
rect 81234 -7654 81854 -2822
rect 84954 50614 85574 86058
rect 88674 198334 89294 222319
rect 88674 198098 88706 198334
rect 88942 198098 89026 198334
rect 89262 198098 89294 198334
rect 88674 198014 89294 198098
rect 88674 197778 88706 198014
rect 88942 197778 89026 198014
rect 89262 197778 89294 198014
rect 88674 162334 89294 197778
rect 88674 162098 88706 162334
rect 88942 162098 89026 162334
rect 89262 162098 89294 162334
rect 88674 162014 89294 162098
rect 88674 161778 88706 162014
rect 88942 161778 89026 162014
rect 89262 161778 89294 162014
rect 88674 126334 89294 161778
rect 88674 126098 88706 126334
rect 88942 126098 89026 126334
rect 89262 126098 89294 126334
rect 88674 126014 89294 126098
rect 88674 125778 88706 126014
rect 88942 125778 89026 126014
rect 89262 125778 89294 126014
rect 88674 90334 89294 125778
rect 92394 202054 93014 222319
rect 92394 201818 92426 202054
rect 92662 201818 92746 202054
rect 92982 201818 93014 202054
rect 92394 201734 93014 201818
rect 92394 201498 92426 201734
rect 92662 201498 92746 201734
rect 92982 201498 93014 201734
rect 92394 166054 93014 201498
rect 92394 165818 92426 166054
rect 92662 165818 92746 166054
rect 92982 165818 93014 166054
rect 92394 165734 93014 165818
rect 92394 165498 92426 165734
rect 92662 165498 92746 165734
rect 92982 165498 93014 165734
rect 92394 130054 93014 165498
rect 92394 129818 92426 130054
rect 92662 129818 92746 130054
rect 92982 129818 93014 130054
rect 92394 129734 93014 129818
rect 92394 129498 92426 129734
rect 92662 129498 92746 129734
rect 92982 129498 93014 129734
rect 92394 111820 93014 129498
rect 96114 205774 96734 241218
rect 96114 205538 96146 205774
rect 96382 205538 96466 205774
rect 96702 205538 96734 205774
rect 96114 205454 96734 205538
rect 96114 205218 96146 205454
rect 96382 205218 96466 205454
rect 96702 205218 96734 205454
rect 96114 169774 96734 205218
rect 96114 169538 96146 169774
rect 96382 169538 96466 169774
rect 96702 169538 96734 169774
rect 96114 169454 96734 169538
rect 96114 169218 96146 169454
rect 96382 169218 96466 169454
rect 96702 169218 96734 169454
rect 96114 133774 96734 169218
rect 96114 133538 96146 133774
rect 96382 133538 96466 133774
rect 96702 133538 96734 133774
rect 96114 133454 96734 133538
rect 96114 133218 96146 133454
rect 96382 133218 96466 133454
rect 96702 133218 96734 133454
rect 96114 111820 96734 133218
rect 99834 711558 100454 711590
rect 99834 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 100454 711558
rect 99834 711238 100454 711322
rect 99834 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 100454 711238
rect 99834 677494 100454 711002
rect 99834 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 100454 677494
rect 99834 677174 100454 677258
rect 99834 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 100454 677174
rect 99834 641494 100454 676938
rect 99834 641258 99866 641494
rect 100102 641258 100186 641494
rect 100422 641258 100454 641494
rect 99834 641174 100454 641258
rect 99834 640938 99866 641174
rect 100102 640938 100186 641174
rect 100422 640938 100454 641174
rect 99834 605494 100454 640938
rect 99834 605258 99866 605494
rect 100102 605258 100186 605494
rect 100422 605258 100454 605494
rect 99834 605174 100454 605258
rect 99834 604938 99866 605174
rect 100102 604938 100186 605174
rect 100422 604938 100454 605174
rect 99834 569494 100454 604938
rect 99834 569258 99866 569494
rect 100102 569258 100186 569494
rect 100422 569258 100454 569494
rect 99834 569174 100454 569258
rect 99834 568938 99866 569174
rect 100102 568938 100186 569174
rect 100422 568938 100454 569174
rect 99834 533494 100454 568938
rect 99834 533258 99866 533494
rect 100102 533258 100186 533494
rect 100422 533258 100454 533494
rect 99834 533174 100454 533258
rect 99834 532938 99866 533174
rect 100102 532938 100186 533174
rect 100422 532938 100454 533174
rect 99834 497494 100454 532938
rect 99834 497258 99866 497494
rect 100102 497258 100186 497494
rect 100422 497258 100454 497494
rect 99834 497174 100454 497258
rect 99834 496938 99866 497174
rect 100102 496938 100186 497174
rect 100422 496938 100454 497174
rect 99834 461494 100454 496938
rect 99834 461258 99866 461494
rect 100102 461258 100186 461494
rect 100422 461258 100454 461494
rect 99834 461174 100454 461258
rect 99834 460938 99866 461174
rect 100102 460938 100186 461174
rect 100422 460938 100454 461174
rect 99834 425494 100454 460938
rect 99834 425258 99866 425494
rect 100102 425258 100186 425494
rect 100422 425258 100454 425494
rect 99834 425174 100454 425258
rect 99834 424938 99866 425174
rect 100102 424938 100186 425174
rect 100422 424938 100454 425174
rect 99834 389494 100454 424938
rect 99834 389258 99866 389494
rect 100102 389258 100186 389494
rect 100422 389258 100454 389494
rect 99834 389174 100454 389258
rect 99834 388938 99866 389174
rect 100102 388938 100186 389174
rect 100422 388938 100454 389174
rect 99834 353494 100454 388938
rect 99834 353258 99866 353494
rect 100102 353258 100186 353494
rect 100422 353258 100454 353494
rect 99834 353174 100454 353258
rect 99834 352938 99866 353174
rect 100102 352938 100186 353174
rect 100422 352938 100454 353174
rect 99834 317494 100454 352938
rect 99834 317258 99866 317494
rect 100102 317258 100186 317494
rect 100422 317258 100454 317494
rect 99834 317174 100454 317258
rect 99834 316938 99866 317174
rect 100102 316938 100186 317174
rect 100422 316938 100454 317174
rect 99834 281494 100454 316938
rect 99834 281258 99866 281494
rect 100102 281258 100186 281494
rect 100422 281258 100454 281494
rect 99834 281174 100454 281258
rect 99834 280938 99866 281174
rect 100102 280938 100186 281174
rect 100422 280938 100454 281174
rect 99834 245494 100454 280938
rect 99834 245258 99866 245494
rect 100102 245258 100186 245494
rect 100422 245258 100454 245494
rect 99834 245174 100454 245258
rect 99834 244938 99866 245174
rect 100102 244938 100186 245174
rect 100422 244938 100454 245174
rect 99834 209494 100454 244938
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 104928 219454 105248 219486
rect 104928 219218 104970 219454
rect 105206 219218 105248 219454
rect 104928 219134 105248 219218
rect 104928 218898 104970 219134
rect 105206 218898 105248 219134
rect 104928 218866 105248 218898
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 99834 209258 99866 209494
rect 100102 209258 100186 209494
rect 100422 209258 100454 209494
rect 99834 209174 100454 209258
rect 99834 208938 99866 209174
rect 100102 208938 100186 209174
rect 100422 208938 100454 209174
rect 99834 173494 100454 208938
rect 99834 173258 99866 173494
rect 100102 173258 100186 173494
rect 100422 173258 100454 173494
rect 99834 173174 100454 173258
rect 99834 172938 99866 173174
rect 100102 172938 100186 173174
rect 100422 172938 100454 173174
rect 99834 137494 100454 172938
rect 99834 137258 99866 137494
rect 100102 137258 100186 137494
rect 100422 137258 100454 137494
rect 99834 137174 100454 137258
rect 99834 136938 99866 137174
rect 100102 136938 100186 137174
rect 100422 136938 100454 137174
rect 99834 111820 100454 136938
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 106043 111212 106109 111213
rect 106043 111210 106044 111212
rect 105678 111150 106044 111210
rect 105678 110941 105738 111150
rect 106043 111148 106044 111150
rect 106108 111148 106109 111212
rect 106043 111147 106109 111148
rect 109794 111134 110414 111218
rect 105675 110940 105741 110941
rect 105675 110876 105676 110940
rect 105740 110876 105741 110940
rect 105675 110875 105741 110876
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 105678 110470 106106 110530
rect 105678 110261 105738 110470
rect 106046 110397 106106 110470
rect 106043 110396 106109 110397
rect 106043 110332 106044 110396
rect 106108 110332 106109 110396
rect 106043 110331 106109 110332
rect 105675 110260 105741 110261
rect 105675 110196 105676 110260
rect 105740 110196 105741 110260
rect 105675 110195 105741 110196
rect 106043 109852 106109 109853
rect 106043 109850 106044 109852
rect 105678 109790 106044 109850
rect 105678 109581 105738 109790
rect 106043 109788 106044 109790
rect 106108 109788 106109 109852
rect 106043 109787 106109 109788
rect 105675 109580 105741 109581
rect 105675 109516 105676 109580
rect 105740 109516 105741 109580
rect 105675 109515 105741 109516
rect 105678 109110 106106 109170
rect 105678 108901 105738 109110
rect 106046 109037 106106 109110
rect 106043 109036 106109 109037
rect 106043 108972 106044 109036
rect 106108 108972 106109 109036
rect 106043 108971 106109 108972
rect 105675 108900 105741 108901
rect 105675 108836 105676 108900
rect 105740 108836 105741 108900
rect 105675 108835 105741 108836
rect 106043 108492 106109 108493
rect 106043 108490 106044 108492
rect 105678 108430 106044 108490
rect 105678 108221 105738 108430
rect 106043 108428 106044 108430
rect 106108 108428 106109 108492
rect 106043 108427 106109 108428
rect 105675 108220 105741 108221
rect 105675 108156 105676 108220
rect 105740 108156 105741 108220
rect 105675 108155 105741 108156
rect 105675 107404 105741 107405
rect 105675 107340 105676 107404
rect 105740 107340 105741 107404
rect 105675 107339 105741 107340
rect 105678 107130 105738 107339
rect 106043 107132 106109 107133
rect 106043 107130 106044 107132
rect 105678 107070 106044 107130
rect 106043 107068 106044 107070
rect 106108 107068 106109 107132
rect 106043 107067 106109 107068
rect 105675 106724 105741 106725
rect 105675 106660 105676 106724
rect 105740 106660 105741 106724
rect 105675 106659 105741 106660
rect 105678 106450 105738 106659
rect 106043 106452 106109 106453
rect 106043 106450 106044 106452
rect 105678 106390 106044 106450
rect 106043 106388 106044 106390
rect 106108 106388 106109 106452
rect 106043 106387 106109 106388
rect 105675 106044 105741 106045
rect 105675 105980 105676 106044
rect 105740 105980 105741 106044
rect 105675 105979 105741 105980
rect 105678 105770 105738 105979
rect 106043 105772 106109 105773
rect 106043 105770 106044 105772
rect 105678 105710 106044 105770
rect 106043 105708 106044 105710
rect 106108 105708 106109 105772
rect 106043 105707 106109 105708
rect 105678 105030 106106 105090
rect 105678 104821 105738 105030
rect 106046 104821 106106 105030
rect 105675 104820 105741 104821
rect 105675 104756 105676 104820
rect 105740 104756 105741 104820
rect 105675 104755 105741 104756
rect 106043 104820 106109 104821
rect 106043 104756 106044 104820
rect 106108 104756 106109 104820
rect 106043 104755 106109 104756
rect 106043 104412 106109 104413
rect 106043 104410 106044 104412
rect 105678 104350 106044 104410
rect 105678 104141 105738 104350
rect 106043 104348 106044 104350
rect 106108 104348 106109 104412
rect 106043 104347 106109 104348
rect 105675 104140 105741 104141
rect 105675 104076 105676 104140
rect 105740 104076 105741 104140
rect 105675 104075 105741 104076
rect 105675 103324 105741 103325
rect 105675 103260 105676 103324
rect 105740 103260 105741 103324
rect 105675 103259 105741 103260
rect 105678 103050 105738 103259
rect 106043 103052 106109 103053
rect 106043 103050 106044 103052
rect 105678 102990 106044 103050
rect 106043 102988 106044 102990
rect 106108 102988 106109 103052
rect 106043 102987 106109 102988
rect 105675 102644 105741 102645
rect 105675 102580 105676 102644
rect 105740 102580 105741 102644
rect 105675 102579 105741 102580
rect 105678 102370 105738 102579
rect 106043 102372 106109 102373
rect 106043 102370 106044 102372
rect 105678 102310 106044 102370
rect 106043 102308 106044 102310
rect 106108 102308 106109 102372
rect 106043 102307 106109 102308
rect 105675 101964 105741 101965
rect 105675 101900 105676 101964
rect 105740 101900 105741 101964
rect 105675 101899 105741 101900
rect 105678 101690 105738 101899
rect 106043 101692 106109 101693
rect 106043 101690 106044 101692
rect 105678 101630 106044 101690
rect 106043 101628 106044 101630
rect 106108 101628 106109 101692
rect 106043 101627 106109 101628
rect 105675 101284 105741 101285
rect 105675 101220 105676 101284
rect 105740 101220 105741 101284
rect 105675 101219 105741 101220
rect 105678 101010 105738 101219
rect 106043 101012 106109 101013
rect 106043 101010 106044 101012
rect 105678 100950 106044 101010
rect 106043 100948 106044 100950
rect 106108 100948 106109 101012
rect 106043 100947 106109 100948
rect 105675 100604 105741 100605
rect 105675 100540 105676 100604
rect 105740 100540 105741 100604
rect 105675 100539 105741 100540
rect 105678 100330 105738 100539
rect 106043 100332 106109 100333
rect 106043 100330 106044 100332
rect 105678 100270 106044 100330
rect 106043 100268 106044 100270
rect 106108 100268 106109 100332
rect 106043 100267 106109 100268
rect 105675 99924 105741 99925
rect 105675 99860 105676 99924
rect 105740 99860 105741 99924
rect 105675 99859 105741 99860
rect 105678 99650 105738 99859
rect 106043 99652 106109 99653
rect 106043 99650 106044 99652
rect 105678 99590 106044 99650
rect 106043 99588 106044 99590
rect 106108 99588 106109 99652
rect 106043 99587 106109 99588
rect 105675 99244 105741 99245
rect 105675 99180 105676 99244
rect 105740 99180 105741 99244
rect 105675 99179 105741 99180
rect 105678 98970 105738 99179
rect 106043 98972 106109 98973
rect 106043 98970 106044 98972
rect 105678 98910 106044 98970
rect 106043 98908 106044 98910
rect 106108 98908 106109 98972
rect 106043 98907 106109 98908
rect 105494 98230 106106 98290
rect 105494 97341 105554 98230
rect 106046 97885 106106 98230
rect 105675 97884 105741 97885
rect 105675 97820 105676 97884
rect 105740 97820 105741 97884
rect 105675 97819 105741 97820
rect 106043 97884 106109 97885
rect 106043 97820 106044 97884
rect 106108 97820 106109 97884
rect 106043 97819 106109 97820
rect 105678 97610 105738 97819
rect 106043 97612 106109 97613
rect 106043 97610 106044 97612
rect 105678 97550 106044 97610
rect 106043 97548 106044 97550
rect 106108 97548 106109 97612
rect 106043 97547 106109 97548
rect 105491 97340 105557 97341
rect 105491 97276 105492 97340
rect 105556 97276 105557 97340
rect 105491 97275 105557 97276
rect 105678 96870 106106 96930
rect 105678 96661 105738 96870
rect 105675 96660 105741 96661
rect 105675 96596 105676 96660
rect 105740 96596 105741 96660
rect 105675 96595 105741 96596
rect 106046 96525 106106 96870
rect 106043 96524 106109 96525
rect 106043 96460 106044 96524
rect 106108 96460 106109 96524
rect 106043 96459 106109 96460
rect 106043 96252 106109 96253
rect 106043 96250 106044 96252
rect 105678 96190 106044 96250
rect 105678 95981 105738 96190
rect 106043 96188 106044 96190
rect 106108 96188 106109 96252
rect 106043 96187 106109 96188
rect 105675 95980 105741 95981
rect 105675 95916 105676 95980
rect 105740 95916 105741 95980
rect 105675 95915 105741 95916
rect 106043 95572 106109 95573
rect 106043 95570 106044 95572
rect 105678 95510 106044 95570
rect 105678 95301 105738 95510
rect 106043 95508 106044 95510
rect 106108 95508 106109 95572
rect 106043 95507 106109 95508
rect 105675 95300 105741 95301
rect 105675 95236 105676 95300
rect 105740 95236 105741 95300
rect 105675 95235 105741 95236
rect 106043 94892 106109 94893
rect 106043 94890 106044 94892
rect 105494 94830 106044 94890
rect 105494 93941 105554 94830
rect 106043 94828 106044 94830
rect 106108 94828 106109 94892
rect 106043 94827 106109 94828
rect 105675 94484 105741 94485
rect 105675 94420 105676 94484
rect 105740 94420 105741 94484
rect 105675 94419 105741 94420
rect 105678 94210 105738 94419
rect 106043 94212 106109 94213
rect 106043 94210 106044 94212
rect 105678 94150 106044 94210
rect 106043 94148 106044 94150
rect 106108 94148 106109 94212
rect 106043 94147 106109 94148
rect 105491 93940 105557 93941
rect 105491 93876 105492 93940
rect 105556 93876 105557 93940
rect 105491 93875 105557 93876
rect 106043 93532 106109 93533
rect 106043 93530 106044 93532
rect 105678 93470 106044 93530
rect 105678 93261 105738 93470
rect 106043 93468 106044 93470
rect 106108 93468 106109 93532
rect 106043 93467 106109 93468
rect 105675 93260 105741 93261
rect 105675 93196 105676 93260
rect 105740 93196 105741 93260
rect 105675 93195 105741 93196
rect 106043 92852 106109 92853
rect 106043 92850 106044 92852
rect 105678 92790 106044 92850
rect 105678 92581 105738 92790
rect 106043 92788 106044 92790
rect 106108 92788 106109 92852
rect 106043 92787 106109 92788
rect 105675 92580 105741 92581
rect 105675 92516 105676 92580
rect 105740 92516 105741 92580
rect 105675 92515 105741 92516
rect 106043 91492 106109 91493
rect 106043 91490 106044 91492
rect 105678 91430 106044 91490
rect 105678 91221 105738 91430
rect 106043 91428 106044 91430
rect 106108 91428 106109 91492
rect 106043 91427 106109 91428
rect 105675 91220 105741 91221
rect 105675 91156 105676 91220
rect 105740 91156 105741 91220
rect 105675 91155 105741 91156
rect 106043 90812 106109 90813
rect 106043 90810 106044 90812
rect 105678 90750 106044 90810
rect 105678 90541 105738 90750
rect 106043 90748 106044 90750
rect 106108 90748 106109 90812
rect 106043 90747 106109 90748
rect 105675 90540 105741 90541
rect 105675 90476 105676 90540
rect 105740 90476 105741 90540
rect 105675 90475 105741 90476
rect 88674 90098 88706 90334
rect 88942 90098 89026 90334
rect 89262 90098 89294 90334
rect 106043 90132 106109 90133
rect 106043 90130 106044 90132
rect 88674 90014 89294 90098
rect 88674 89778 88706 90014
rect 88942 89778 89026 90014
rect 89262 89778 89294 90014
rect 105678 90070 106044 90130
rect 105678 89861 105738 90070
rect 106043 90068 106044 90070
rect 106108 90068 106109 90132
rect 106043 90067 106109 90068
rect 105675 89860 105741 89861
rect 105675 89796 105676 89860
rect 105740 89796 105741 89860
rect 105675 89795 105741 89796
rect 87825 79174 88145 79206
rect 87825 78938 87867 79174
rect 88103 78938 88145 79174
rect 87825 78854 88145 78938
rect 87825 78618 87867 78854
rect 88103 78618 88145 78854
rect 87825 78586 88145 78618
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 84954 -3226 85574 14058
rect 84954 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 85574 -3226
rect 84954 -3546 85574 -3462
rect 84954 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 85574 -3546
rect 84954 -7654 85574 -3782
rect 88674 54334 89294 89778
rect 106043 89452 106109 89453
rect 106043 89450 106044 89452
rect 105678 89390 106044 89450
rect 105678 89181 105738 89390
rect 106043 89388 106044 89390
rect 106108 89388 106109 89452
rect 106043 89387 106109 89388
rect 105675 89180 105741 89181
rect 105675 89116 105676 89180
rect 105740 89116 105741 89180
rect 105675 89115 105741 89116
rect 106043 88772 106109 88773
rect 106043 88770 106044 88772
rect 105678 88710 106044 88770
rect 105678 88501 105738 88710
rect 106043 88708 106044 88710
rect 106108 88708 106109 88772
rect 106043 88707 106109 88708
rect 105675 88500 105741 88501
rect 105675 88436 105676 88500
rect 105740 88436 105741 88500
rect 105675 88435 105741 88436
rect 106043 88092 106109 88093
rect 106043 88090 106044 88092
rect 105678 88030 106044 88090
rect 105678 87821 105738 88030
rect 106043 88028 106044 88030
rect 106108 88028 106109 88092
rect 106043 88027 106109 88028
rect 105675 87820 105741 87821
rect 105675 87756 105676 87820
rect 105740 87756 105741 87820
rect 105675 87755 105741 87756
rect 106043 87412 106109 87413
rect 106043 87410 106044 87412
rect 105678 87350 106044 87410
rect 105678 87141 105738 87350
rect 106043 87348 106044 87350
rect 106108 87348 106109 87412
rect 106043 87347 106109 87348
rect 105675 87140 105741 87141
rect 105675 87076 105676 87140
rect 105740 87076 105741 87140
rect 105675 87075 105741 87076
rect 106043 86732 106109 86733
rect 106043 86730 106044 86732
rect 105678 86670 106044 86730
rect 105678 86461 105738 86670
rect 106043 86668 106044 86670
rect 106108 86668 106109 86732
rect 106043 86667 106109 86668
rect 105675 86460 105741 86461
rect 105675 86396 105676 86460
rect 105740 86396 105741 86460
rect 105675 86395 105741 86396
rect 106043 86052 106109 86053
rect 106043 86050 106044 86052
rect 105678 85990 106044 86050
rect 105678 85781 105738 85990
rect 106043 85988 106044 85990
rect 106108 85988 106109 86052
rect 106043 85987 106109 85988
rect 105675 85780 105741 85781
rect 105675 85716 105676 85780
rect 105740 85716 105741 85780
rect 105675 85715 105741 85716
rect 106043 84692 106109 84693
rect 106043 84690 106044 84692
rect 105678 84630 106044 84690
rect 105678 84421 105738 84630
rect 106043 84628 106044 84630
rect 106108 84628 106109 84692
rect 106043 84627 106109 84628
rect 105675 84420 105741 84421
rect 105675 84356 105676 84420
rect 105740 84356 105741 84420
rect 105675 84355 105741 84356
rect 106043 84012 106109 84013
rect 106043 84010 106044 84012
rect 105678 83950 106044 84010
rect 105678 83741 105738 83950
rect 106043 83948 106044 83950
rect 106108 83948 106109 84012
rect 106043 83947 106109 83948
rect 105675 83740 105741 83741
rect 105675 83676 105676 83740
rect 105740 83676 105741 83740
rect 105675 83675 105741 83676
rect 106043 83332 106109 83333
rect 106043 83330 106044 83332
rect 105678 83270 106044 83330
rect 105678 83061 105738 83270
rect 106043 83268 106044 83270
rect 106108 83268 106109 83332
rect 106043 83267 106109 83268
rect 106779 83196 106845 83197
rect 106779 83132 106780 83196
rect 106844 83132 106845 83196
rect 106779 83131 106845 83132
rect 105675 83060 105741 83061
rect 105675 82996 105676 83060
rect 105740 82996 105741 83060
rect 105675 82995 105741 82996
rect 106043 82652 106109 82653
rect 106043 82650 106044 82652
rect 105678 82590 106044 82650
rect 105678 82381 105738 82590
rect 106043 82588 106044 82590
rect 106108 82588 106109 82652
rect 106043 82587 106109 82588
rect 105675 82380 105741 82381
rect 105675 82316 105676 82380
rect 105740 82316 105741 82380
rect 105675 82315 105741 82316
rect 106043 81972 106109 81973
rect 106043 81970 106044 81972
rect 105678 81910 106044 81970
rect 105678 81701 105738 81910
rect 106043 81908 106044 81910
rect 106108 81908 106109 81972
rect 106043 81907 106109 81908
rect 106227 81836 106293 81837
rect 106227 81772 106228 81836
rect 106292 81772 106293 81836
rect 106227 81771 106293 81772
rect 105675 81700 105741 81701
rect 105675 81636 105676 81700
rect 105740 81636 105741 81700
rect 105675 81635 105741 81636
rect 106043 81292 106109 81293
rect 106043 81290 106044 81292
rect 105678 81230 106044 81290
rect 105678 81021 105738 81230
rect 106043 81228 106044 81230
rect 106108 81228 106109 81292
rect 106043 81227 106109 81228
rect 105675 81020 105741 81021
rect 105675 80956 105676 81020
rect 105740 80956 105741 81020
rect 105675 80955 105741 80956
rect 106043 80612 106109 80613
rect 106043 80610 106044 80612
rect 105678 80550 106044 80610
rect 105678 80341 105738 80550
rect 106043 80548 106044 80550
rect 106108 80548 106109 80612
rect 106043 80547 106109 80548
rect 105675 80340 105741 80341
rect 105675 80276 105676 80340
rect 105740 80276 105741 80340
rect 105675 80275 105741 80276
rect 106230 80070 106290 81771
rect 105310 80010 106290 80070
rect 96266 79174 96586 79206
rect 96266 78938 96308 79174
rect 96544 78938 96586 79174
rect 96266 78854 96586 78938
rect 96266 78618 96308 78854
rect 96544 78618 96586 78854
rect 96266 78586 96586 78618
rect 104707 79174 105027 79206
rect 104707 78938 104749 79174
rect 104985 78938 105027 79174
rect 104707 78854 105027 78938
rect 104707 78618 104749 78854
rect 104985 78618 105027 78854
rect 104707 78586 105027 78618
rect 105310 77310 105370 80010
rect 106043 79932 106109 79933
rect 106043 79930 106044 79932
rect 105678 79870 106044 79930
rect 105678 79661 105738 79870
rect 106043 79868 106044 79870
rect 106108 79868 106109 79932
rect 106043 79867 106109 79868
rect 105675 79660 105741 79661
rect 105675 79596 105676 79660
rect 105740 79596 105741 79660
rect 105675 79595 105741 79596
rect 106043 79252 106109 79253
rect 106043 79250 106044 79252
rect 105678 79190 106044 79250
rect 105678 78981 105738 79190
rect 106043 79188 106044 79190
rect 106108 79188 106109 79252
rect 106043 79187 106109 79188
rect 105675 78980 105741 78981
rect 105675 78916 105676 78980
rect 105740 78916 105741 78980
rect 105675 78915 105741 78916
rect 106043 77892 106109 77893
rect 106043 77890 106044 77892
rect 105678 77830 106044 77890
rect 105678 77621 105738 77830
rect 106043 77828 106044 77830
rect 106108 77828 106109 77892
rect 106043 77827 106109 77828
rect 105675 77620 105741 77621
rect 105675 77556 105676 77620
rect 105740 77556 105741 77620
rect 105675 77555 105741 77556
rect 105126 77250 105370 77310
rect 92046 75454 92366 75486
rect 92046 75218 92088 75454
rect 92324 75218 92366 75454
rect 92046 75134 92366 75218
rect 92046 74898 92088 75134
rect 92324 74898 92366 75134
rect 92046 74866 92366 74898
rect 100487 75454 100807 75486
rect 100487 75218 100529 75454
rect 100765 75218 100807 75454
rect 100487 75134 100807 75218
rect 100487 74898 100529 75134
rect 100765 74898 100807 75134
rect 100487 74866 100807 74898
rect 105126 74490 105186 77250
rect 105675 76804 105741 76805
rect 105675 76740 105676 76804
rect 105740 76740 105741 76804
rect 105675 76739 105741 76740
rect 105678 76530 105738 76739
rect 106043 76532 106109 76533
rect 106043 76530 106044 76532
rect 105678 76470 106044 76530
rect 106043 76468 106044 76470
rect 106108 76468 106109 76532
rect 106043 76467 106109 76468
rect 106411 76532 106477 76533
rect 106411 76468 106412 76532
rect 106476 76468 106477 76532
rect 106411 76467 106477 76468
rect 105675 76124 105741 76125
rect 105675 76060 105676 76124
rect 105740 76060 105741 76124
rect 105675 76059 105741 76060
rect 105678 75850 105738 76059
rect 106043 75988 106109 75989
rect 106043 75924 106044 75988
rect 106108 75924 106109 75988
rect 106043 75923 106109 75924
rect 106046 75850 106106 75923
rect 105678 75790 106106 75850
rect 106043 75716 106109 75717
rect 106043 75652 106044 75716
rect 106108 75652 106109 75716
rect 106043 75651 106109 75652
rect 105675 75580 105741 75581
rect 105675 75516 105676 75580
rect 105740 75578 105741 75580
rect 106046 75578 106106 75651
rect 105740 75518 106106 75578
rect 105740 75516 105741 75518
rect 105675 75515 105741 75516
rect 106043 75172 106109 75173
rect 106043 75108 106044 75172
rect 106108 75108 106109 75172
rect 106414 75170 106474 76467
rect 106043 75107 106109 75108
rect 106230 75110 106474 75170
rect 105675 74900 105741 74901
rect 105675 74836 105676 74900
rect 105740 74898 105741 74900
rect 106046 74898 106106 75107
rect 106230 75037 106290 75110
rect 106227 75036 106293 75037
rect 106227 74972 106228 75036
rect 106292 74972 106293 75036
rect 106227 74971 106293 74972
rect 105740 74838 106106 74898
rect 105740 74836 105741 74838
rect 105675 74835 105741 74836
rect 105126 74430 105370 74490
rect 88674 54098 88706 54334
rect 88942 54098 89026 54334
rect 89262 54098 89294 54334
rect 88674 54014 89294 54098
rect 88674 53778 88706 54014
rect 88942 53778 89026 54014
rect 89262 53778 89294 54014
rect 88674 18334 89294 53778
rect 88674 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 89294 18334
rect 88674 18014 89294 18098
rect 88674 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 89294 18014
rect 88674 -4186 89294 17778
rect 88674 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 89294 -4186
rect 88674 -4506 89294 -4422
rect 88674 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 89294 -4506
rect 88674 -7654 89294 -4742
rect 92394 58054 93014 70068
rect 92394 57818 92426 58054
rect 92662 57818 92746 58054
rect 92982 57818 93014 58054
rect 92394 57734 93014 57818
rect 92394 57498 92426 57734
rect 92662 57498 92746 57734
rect 92982 57498 93014 57734
rect 92394 22054 93014 57498
rect 92394 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 93014 22054
rect 92394 21734 93014 21818
rect 92394 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 93014 21734
rect 92394 -5146 93014 21498
rect 92394 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 93014 -5146
rect 92394 -5466 93014 -5382
rect 92394 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 93014 -5466
rect 92394 -7654 93014 -5702
rect 96114 61774 96734 70068
rect 96114 61538 96146 61774
rect 96382 61538 96466 61774
rect 96702 61538 96734 61774
rect 96114 61454 96734 61538
rect 96114 61218 96146 61454
rect 96382 61218 96466 61454
rect 96702 61218 96734 61454
rect 96114 25774 96734 61218
rect 96114 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 96734 25774
rect 96114 25454 96734 25538
rect 96114 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 96734 25454
rect 96114 -6106 96734 25218
rect 96114 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 96734 -6106
rect 96114 -6426 96734 -6342
rect 96114 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 96734 -6426
rect 96114 -7654 96734 -6662
rect 99834 65494 100454 70068
rect 105310 67285 105370 74430
rect 105675 74084 105741 74085
rect 105675 74020 105676 74084
rect 105740 74020 105741 74084
rect 105675 74019 105741 74020
rect 106043 74084 106109 74085
rect 106043 74020 106044 74084
rect 106108 74020 106109 74084
rect 106043 74019 106109 74020
rect 105678 73810 105738 74019
rect 106046 73810 106106 74019
rect 105678 73750 106106 73810
rect 106043 73676 106109 73677
rect 106043 73612 106044 73676
rect 106108 73612 106109 73676
rect 106043 73611 106109 73612
rect 106046 73538 106106 73611
rect 105678 73478 106106 73538
rect 105678 73405 105738 73478
rect 105675 73404 105741 73405
rect 105675 73340 105676 73404
rect 105740 73340 105741 73404
rect 105675 73339 105741 73340
rect 106043 72860 106109 72861
rect 106043 72796 106044 72860
rect 106108 72796 106109 72860
rect 106043 72795 106109 72796
rect 105675 72724 105741 72725
rect 105675 72660 105676 72724
rect 105740 72660 105741 72724
rect 105675 72659 105741 72660
rect 105678 72450 105738 72659
rect 106046 72450 106106 72795
rect 105678 72390 106106 72450
rect 106043 72316 106109 72317
rect 106043 72252 106044 72316
rect 106108 72252 106109 72316
rect 106043 72251 106109 72252
rect 105675 72180 105741 72181
rect 105675 72116 105676 72180
rect 105740 72178 105741 72180
rect 106046 72178 106106 72251
rect 105740 72118 106106 72178
rect 105740 72116 105741 72118
rect 105675 72115 105741 72116
rect 106043 71092 106109 71093
rect 106043 71028 106044 71092
rect 106108 71028 106109 71092
rect 106043 71027 106109 71028
rect 105675 70684 105741 70685
rect 105675 70620 105676 70684
rect 105740 70620 105741 70684
rect 105675 70619 105741 70620
rect 105678 70410 105738 70619
rect 106046 70410 106106 71027
rect 105494 70350 105738 70410
rect 105862 70350 106106 70410
rect 105494 69325 105554 70350
rect 105675 70140 105741 70141
rect 105675 70076 105676 70140
rect 105740 70076 105741 70140
rect 105675 70075 105741 70076
rect 105678 69730 105738 70075
rect 105862 69730 105922 70350
rect 106043 70276 106109 70277
rect 106043 70212 106044 70276
rect 106108 70212 106109 70276
rect 106043 70211 106109 70212
rect 105678 69670 105922 69730
rect 106046 69461 106106 70211
rect 106782 69597 106842 83131
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 106779 69596 106845 69597
rect 106779 69532 106780 69596
rect 106844 69532 106845 69596
rect 106779 69531 106845 69532
rect 106043 69460 106109 69461
rect 106043 69396 106044 69460
rect 106108 69396 106109 69460
rect 106043 69395 106109 69396
rect 105491 69324 105557 69325
rect 105491 69260 105492 69324
rect 105556 69260 105557 69324
rect 105491 69259 105557 69260
rect 105307 67284 105373 67285
rect 105307 67220 105308 67284
rect 105372 67220 105373 67284
rect 105307 67219 105373 67220
rect 99834 65258 99866 65494
rect 100102 65258 100186 65494
rect 100422 65258 100454 65494
rect 99834 65174 100454 65258
rect 99834 64938 99866 65174
rect 100102 64938 100186 65174
rect 100422 64938 100454 65174
rect 99834 29494 100454 64938
rect 99834 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 100454 29494
rect 99834 29174 100454 29258
rect 99834 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 100454 29174
rect 99834 -7066 100454 28938
rect 99834 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 100454 -7066
rect 99834 -7386 100454 -7302
rect 99834 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 100454 -7386
rect 99834 -7654 100454 -7622
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 113514 705798 114134 711590
rect 113514 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 114134 705798
rect 113514 705478 114134 705562
rect 113514 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 114134 705478
rect 113514 691174 114134 705242
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -1306 114134 6618
rect 113514 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 114134 -1306
rect 113514 -1626 114134 -1542
rect 113514 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 114134 -1626
rect 113514 -7654 114134 -1862
rect 117234 706758 117854 711590
rect 117234 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 117854 706758
rect 117234 706438 117854 706522
rect 117234 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 117854 706438
rect 117234 694894 117854 706202
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 120954 707718 121574 711590
rect 120954 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 121574 707718
rect 120954 707398 121574 707482
rect 120954 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 121574 707398
rect 120954 698614 121574 707162
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120027 251972 120093 251973
rect 120027 251908 120028 251972
rect 120092 251908 120093 251972
rect 120027 251907 120093 251908
rect 119843 251564 119909 251565
rect 119843 251500 119844 251564
rect 119908 251500 119909 251564
rect 119843 251499 119909 251500
rect 119475 250204 119541 250205
rect 119475 250140 119476 250204
rect 119540 250140 119541 250204
rect 119475 250139 119541 250140
rect 119478 232525 119538 250139
rect 119659 250068 119725 250069
rect 119659 250004 119660 250068
rect 119724 250004 119725 250068
rect 119659 250003 119725 250004
rect 119662 238770 119722 250003
rect 119846 248029 119906 251499
rect 119843 248028 119909 248029
rect 119843 247964 119844 248028
rect 119908 247964 119909 248028
rect 119843 247963 119909 247964
rect 120030 247621 120090 251907
rect 120027 247620 120093 247621
rect 120027 247556 120028 247620
rect 120092 247556 120093 247620
rect 120027 247555 120093 247556
rect 120211 240276 120277 240277
rect 120211 240212 120212 240276
rect 120276 240212 120277 240276
rect 120211 240211 120277 240212
rect 119662 238710 119906 238770
rect 119846 233069 119906 238710
rect 119843 233068 119909 233069
rect 119843 233004 119844 233068
rect 119908 233004 119909 233068
rect 119843 233003 119909 233004
rect 119475 232524 119541 232525
rect 119475 232460 119476 232524
rect 119540 232460 119541 232524
rect 119475 232459 119541 232460
rect 119659 229260 119725 229261
rect 119659 229196 119660 229260
rect 119724 229196 119725 229260
rect 119659 229195 119725 229196
rect 119291 228580 119357 228581
rect 119291 228516 119292 228580
rect 119356 228516 119357 228580
rect 119291 228515 119357 228516
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 119294 225450 119354 228515
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 118926 225390 119354 225450
rect 118926 125357 118986 225390
rect 119291 221236 119357 221237
rect 119291 221172 119292 221236
rect 119356 221172 119357 221236
rect 119291 221171 119357 221172
rect 119294 219450 119354 221171
rect 119110 219390 119354 219450
rect 119110 165613 119170 219390
rect 119291 210764 119357 210765
rect 119291 210700 119292 210764
rect 119356 210700 119357 210764
rect 119291 210699 119357 210700
rect 119294 196757 119354 210699
rect 119291 196756 119357 196757
rect 119291 196692 119292 196756
rect 119356 196692 119357 196756
rect 119291 196691 119357 196692
rect 119107 165612 119173 165613
rect 119107 165548 119108 165612
rect 119172 165548 119173 165612
rect 119107 165547 119173 165548
rect 119662 125493 119722 229195
rect 120027 227900 120093 227901
rect 120027 227836 120028 227900
rect 120092 227836 120093 227900
rect 120027 227835 120093 227836
rect 119659 125492 119725 125493
rect 119659 125428 119660 125492
rect 119724 125428 119725 125492
rect 119659 125427 119725 125428
rect 118923 125356 118989 125357
rect 118923 125292 118924 125356
rect 118988 125292 118989 125356
rect 118923 125291 118989 125292
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 120030 95301 120090 227835
rect 120214 196621 120274 240211
rect 120954 230614 121574 266058
rect 124674 708678 125294 711590
rect 124674 708442 124706 708678
rect 124942 708442 125026 708678
rect 125262 708442 125294 708678
rect 124674 708358 125294 708442
rect 124674 708122 124706 708358
rect 124942 708122 125026 708358
rect 125262 708122 125294 708358
rect 124674 666334 125294 708122
rect 124674 666098 124706 666334
rect 124942 666098 125026 666334
rect 125262 666098 125294 666334
rect 124674 666014 125294 666098
rect 124674 665778 124706 666014
rect 124942 665778 125026 666014
rect 125262 665778 125294 666014
rect 124674 630334 125294 665778
rect 124674 630098 124706 630334
rect 124942 630098 125026 630334
rect 125262 630098 125294 630334
rect 124674 630014 125294 630098
rect 124674 629778 124706 630014
rect 124942 629778 125026 630014
rect 125262 629778 125294 630014
rect 124674 594334 125294 629778
rect 124674 594098 124706 594334
rect 124942 594098 125026 594334
rect 125262 594098 125294 594334
rect 124674 594014 125294 594098
rect 124674 593778 124706 594014
rect 124942 593778 125026 594014
rect 125262 593778 125294 594014
rect 124674 558334 125294 593778
rect 124674 558098 124706 558334
rect 124942 558098 125026 558334
rect 125262 558098 125294 558334
rect 124674 558014 125294 558098
rect 124674 557778 124706 558014
rect 124942 557778 125026 558014
rect 125262 557778 125294 558014
rect 124674 522334 125294 557778
rect 124674 522098 124706 522334
rect 124942 522098 125026 522334
rect 125262 522098 125294 522334
rect 124674 522014 125294 522098
rect 124674 521778 124706 522014
rect 124942 521778 125026 522014
rect 125262 521778 125294 522014
rect 124674 486334 125294 521778
rect 124674 486098 124706 486334
rect 124942 486098 125026 486334
rect 125262 486098 125294 486334
rect 124674 486014 125294 486098
rect 124674 485778 124706 486014
rect 124942 485778 125026 486014
rect 125262 485778 125294 486014
rect 124674 450334 125294 485778
rect 124674 450098 124706 450334
rect 124942 450098 125026 450334
rect 125262 450098 125294 450334
rect 124674 450014 125294 450098
rect 124674 449778 124706 450014
rect 124942 449778 125026 450014
rect 125262 449778 125294 450014
rect 124674 414334 125294 449778
rect 124674 414098 124706 414334
rect 124942 414098 125026 414334
rect 125262 414098 125294 414334
rect 124674 414014 125294 414098
rect 124674 413778 124706 414014
rect 124942 413778 125026 414014
rect 125262 413778 125294 414014
rect 124674 378334 125294 413778
rect 124674 378098 124706 378334
rect 124942 378098 125026 378334
rect 125262 378098 125294 378334
rect 124674 378014 125294 378098
rect 124674 377778 124706 378014
rect 124942 377778 125026 378014
rect 125262 377778 125294 378014
rect 124674 342334 125294 377778
rect 124674 342098 124706 342334
rect 124942 342098 125026 342334
rect 125262 342098 125294 342334
rect 124674 342014 125294 342098
rect 124674 341778 124706 342014
rect 124942 341778 125026 342014
rect 125262 341778 125294 342014
rect 124674 306334 125294 341778
rect 124674 306098 124706 306334
rect 124942 306098 125026 306334
rect 125262 306098 125294 306334
rect 124674 306014 125294 306098
rect 124674 305778 124706 306014
rect 124942 305778 125026 306014
rect 125262 305778 125294 306014
rect 124674 270334 125294 305778
rect 124674 270098 124706 270334
rect 124942 270098 125026 270334
rect 125262 270098 125294 270334
rect 124674 270014 125294 270098
rect 124674 269778 124706 270014
rect 124942 269778 125026 270014
rect 125262 269778 125294 270014
rect 121867 246260 121933 246261
rect 121867 246196 121868 246260
rect 121932 246196 121933 246260
rect 121867 246195 121933 246196
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120579 226404 120645 226405
rect 120579 226340 120580 226404
rect 120644 226340 120645 226404
rect 120579 226339 120645 226340
rect 120211 196620 120277 196621
rect 120211 196556 120212 196620
rect 120276 196556 120277 196620
rect 120211 196555 120277 196556
rect 120582 166973 120642 226339
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120579 166972 120645 166973
rect 120579 166908 120580 166972
rect 120644 166908 120645 166972
rect 120579 166907 120645 166908
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 121870 123453 121930 246195
rect 122235 242996 122301 242997
rect 122235 242932 122236 242996
rect 122300 242932 122301 242996
rect 122235 242931 122301 242932
rect 122051 213076 122117 213077
rect 122051 213012 122052 213076
rect 122116 213012 122117 213076
rect 122051 213011 122117 213012
rect 121867 123452 121933 123453
rect 121867 123388 121868 123452
rect 121932 123388 121933 123452
rect 121867 123387 121933 123388
rect 122054 122909 122114 213011
rect 122238 192541 122298 242931
rect 124674 234334 125294 269778
rect 124674 234098 124706 234334
rect 124942 234098 125026 234334
rect 125262 234098 125294 234334
rect 124674 234014 125294 234098
rect 124674 233778 124706 234014
rect 124942 233778 125026 234014
rect 125262 233778 125294 234014
rect 122419 210220 122485 210221
rect 122419 210156 122420 210220
rect 122484 210156 122485 210220
rect 122419 210155 122485 210156
rect 122235 192540 122301 192541
rect 122235 192476 122236 192540
rect 122300 192476 122301 192540
rect 122235 192475 122301 192476
rect 122422 175949 122482 210155
rect 124674 198334 125294 233778
rect 124674 198098 124706 198334
rect 124942 198098 125026 198334
rect 125262 198098 125294 198334
rect 124674 198014 125294 198098
rect 124674 197778 124706 198014
rect 124942 197778 125026 198014
rect 125262 197778 125294 198014
rect 122419 175948 122485 175949
rect 122419 175884 122420 175948
rect 122484 175884 122485 175948
rect 122419 175883 122485 175884
rect 124674 162334 125294 197778
rect 124674 162098 124706 162334
rect 124942 162098 125026 162334
rect 125262 162098 125294 162334
rect 124674 162014 125294 162098
rect 124674 161778 124706 162014
rect 124942 161778 125026 162014
rect 125262 161778 125294 162014
rect 124674 126334 125294 161778
rect 124674 126098 124706 126334
rect 124942 126098 125026 126334
rect 125262 126098 125294 126334
rect 124674 126014 125294 126098
rect 124674 125778 124706 126014
rect 124942 125778 125026 126014
rect 125262 125778 125294 126014
rect 122051 122908 122117 122909
rect 122051 122844 122052 122908
rect 122116 122844 122117 122908
rect 122051 122843 122117 122844
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120027 95300 120093 95301
rect 120027 95236 120028 95300
rect 120092 95236 120093 95300
rect 120027 95235 120093 95236
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -2266 117854 10338
rect 117234 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 117854 -2266
rect 117234 -2586 117854 -2502
rect 117234 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 117854 -2586
rect 117234 -7654 117854 -2822
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 120954 -3226 121574 14058
rect 120954 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 121574 -3226
rect 120954 -3546 121574 -3462
rect 120954 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 121574 -3546
rect 120954 -7654 121574 -3782
rect 124674 90334 125294 125778
rect 124674 90098 124706 90334
rect 124942 90098 125026 90334
rect 125262 90098 125294 90334
rect 124674 90014 125294 90098
rect 124674 89778 124706 90014
rect 124942 89778 125026 90014
rect 125262 89778 125294 90014
rect 124674 54334 125294 89778
rect 124674 54098 124706 54334
rect 124942 54098 125026 54334
rect 125262 54098 125294 54334
rect 124674 54014 125294 54098
rect 124674 53778 124706 54014
rect 124942 53778 125026 54014
rect 125262 53778 125294 54014
rect 124674 18334 125294 53778
rect 124674 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 125294 18334
rect 124674 18014 125294 18098
rect 124674 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 125294 18014
rect 124674 -4186 125294 17778
rect 124674 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 125294 -4186
rect 124674 -4506 125294 -4422
rect 124674 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 125294 -4506
rect 124674 -7654 125294 -4742
rect 128394 709638 129014 711590
rect 128394 709402 128426 709638
rect 128662 709402 128746 709638
rect 128982 709402 129014 709638
rect 128394 709318 129014 709402
rect 128394 709082 128426 709318
rect 128662 709082 128746 709318
rect 128982 709082 129014 709318
rect 128394 670054 129014 709082
rect 128394 669818 128426 670054
rect 128662 669818 128746 670054
rect 128982 669818 129014 670054
rect 128394 669734 129014 669818
rect 128394 669498 128426 669734
rect 128662 669498 128746 669734
rect 128982 669498 129014 669734
rect 128394 634054 129014 669498
rect 128394 633818 128426 634054
rect 128662 633818 128746 634054
rect 128982 633818 129014 634054
rect 128394 633734 129014 633818
rect 128394 633498 128426 633734
rect 128662 633498 128746 633734
rect 128982 633498 129014 633734
rect 128394 598054 129014 633498
rect 128394 597818 128426 598054
rect 128662 597818 128746 598054
rect 128982 597818 129014 598054
rect 128394 597734 129014 597818
rect 128394 597498 128426 597734
rect 128662 597498 128746 597734
rect 128982 597498 129014 597734
rect 128394 562054 129014 597498
rect 128394 561818 128426 562054
rect 128662 561818 128746 562054
rect 128982 561818 129014 562054
rect 128394 561734 129014 561818
rect 128394 561498 128426 561734
rect 128662 561498 128746 561734
rect 128982 561498 129014 561734
rect 128394 526054 129014 561498
rect 128394 525818 128426 526054
rect 128662 525818 128746 526054
rect 128982 525818 129014 526054
rect 128394 525734 129014 525818
rect 128394 525498 128426 525734
rect 128662 525498 128746 525734
rect 128982 525498 129014 525734
rect 128394 490054 129014 525498
rect 128394 489818 128426 490054
rect 128662 489818 128746 490054
rect 128982 489818 129014 490054
rect 128394 489734 129014 489818
rect 128394 489498 128426 489734
rect 128662 489498 128746 489734
rect 128982 489498 129014 489734
rect 128394 454054 129014 489498
rect 128394 453818 128426 454054
rect 128662 453818 128746 454054
rect 128982 453818 129014 454054
rect 128394 453734 129014 453818
rect 128394 453498 128426 453734
rect 128662 453498 128746 453734
rect 128982 453498 129014 453734
rect 128394 418054 129014 453498
rect 128394 417818 128426 418054
rect 128662 417818 128746 418054
rect 128982 417818 129014 418054
rect 128394 417734 129014 417818
rect 128394 417498 128426 417734
rect 128662 417498 128746 417734
rect 128982 417498 129014 417734
rect 128394 382054 129014 417498
rect 128394 381818 128426 382054
rect 128662 381818 128746 382054
rect 128982 381818 129014 382054
rect 128394 381734 129014 381818
rect 128394 381498 128426 381734
rect 128662 381498 128746 381734
rect 128982 381498 129014 381734
rect 128394 346054 129014 381498
rect 128394 345818 128426 346054
rect 128662 345818 128746 346054
rect 128982 345818 129014 346054
rect 128394 345734 129014 345818
rect 128394 345498 128426 345734
rect 128662 345498 128746 345734
rect 128982 345498 129014 345734
rect 128394 310054 129014 345498
rect 128394 309818 128426 310054
rect 128662 309818 128746 310054
rect 128982 309818 129014 310054
rect 128394 309734 129014 309818
rect 128394 309498 128426 309734
rect 128662 309498 128746 309734
rect 128982 309498 129014 309734
rect 128394 274054 129014 309498
rect 128394 273818 128426 274054
rect 128662 273818 128746 274054
rect 128982 273818 129014 274054
rect 128394 273734 129014 273818
rect 128394 273498 128426 273734
rect 128662 273498 128746 273734
rect 128982 273498 129014 273734
rect 128394 238054 129014 273498
rect 128394 237818 128426 238054
rect 128662 237818 128746 238054
rect 128982 237818 129014 238054
rect 128394 237734 129014 237818
rect 128394 237498 128426 237734
rect 128662 237498 128746 237734
rect 128982 237498 129014 237734
rect 128394 202054 129014 237498
rect 128394 201818 128426 202054
rect 128662 201818 128746 202054
rect 128982 201818 129014 202054
rect 128394 201734 129014 201818
rect 128394 201498 128426 201734
rect 128662 201498 128746 201734
rect 128982 201498 129014 201734
rect 128394 166054 129014 201498
rect 128394 165818 128426 166054
rect 128662 165818 128746 166054
rect 128982 165818 129014 166054
rect 128394 165734 129014 165818
rect 128394 165498 128426 165734
rect 128662 165498 128746 165734
rect 128982 165498 129014 165734
rect 128394 130054 129014 165498
rect 128394 129818 128426 130054
rect 128662 129818 128746 130054
rect 128982 129818 129014 130054
rect 128394 129734 129014 129818
rect 128394 129498 128426 129734
rect 128662 129498 128746 129734
rect 128982 129498 129014 129734
rect 128394 94054 129014 129498
rect 128394 93818 128426 94054
rect 128662 93818 128746 94054
rect 128982 93818 129014 94054
rect 128394 93734 129014 93818
rect 128394 93498 128426 93734
rect 128662 93498 128746 93734
rect 128982 93498 129014 93734
rect 128394 58054 129014 93498
rect 128394 57818 128426 58054
rect 128662 57818 128746 58054
rect 128982 57818 129014 58054
rect 128394 57734 129014 57818
rect 128394 57498 128426 57734
rect 128662 57498 128746 57734
rect 128982 57498 129014 57734
rect 128394 22054 129014 57498
rect 128394 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 129014 22054
rect 128394 21734 129014 21818
rect 128394 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 129014 21734
rect 128394 -5146 129014 21498
rect 128394 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 129014 -5146
rect 128394 -5466 129014 -5382
rect 128394 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 129014 -5466
rect 128394 -7654 129014 -5702
rect 132114 710598 132734 711590
rect 132114 710362 132146 710598
rect 132382 710362 132466 710598
rect 132702 710362 132734 710598
rect 132114 710278 132734 710362
rect 132114 710042 132146 710278
rect 132382 710042 132466 710278
rect 132702 710042 132734 710278
rect 132114 673774 132734 710042
rect 132114 673538 132146 673774
rect 132382 673538 132466 673774
rect 132702 673538 132734 673774
rect 132114 673454 132734 673538
rect 132114 673218 132146 673454
rect 132382 673218 132466 673454
rect 132702 673218 132734 673454
rect 132114 637774 132734 673218
rect 132114 637538 132146 637774
rect 132382 637538 132466 637774
rect 132702 637538 132734 637774
rect 132114 637454 132734 637538
rect 132114 637218 132146 637454
rect 132382 637218 132466 637454
rect 132702 637218 132734 637454
rect 132114 601774 132734 637218
rect 132114 601538 132146 601774
rect 132382 601538 132466 601774
rect 132702 601538 132734 601774
rect 132114 601454 132734 601538
rect 132114 601218 132146 601454
rect 132382 601218 132466 601454
rect 132702 601218 132734 601454
rect 132114 565774 132734 601218
rect 132114 565538 132146 565774
rect 132382 565538 132466 565774
rect 132702 565538 132734 565774
rect 132114 565454 132734 565538
rect 132114 565218 132146 565454
rect 132382 565218 132466 565454
rect 132702 565218 132734 565454
rect 132114 529774 132734 565218
rect 132114 529538 132146 529774
rect 132382 529538 132466 529774
rect 132702 529538 132734 529774
rect 132114 529454 132734 529538
rect 132114 529218 132146 529454
rect 132382 529218 132466 529454
rect 132702 529218 132734 529454
rect 132114 493774 132734 529218
rect 132114 493538 132146 493774
rect 132382 493538 132466 493774
rect 132702 493538 132734 493774
rect 132114 493454 132734 493538
rect 132114 493218 132146 493454
rect 132382 493218 132466 493454
rect 132702 493218 132734 493454
rect 132114 457774 132734 493218
rect 132114 457538 132146 457774
rect 132382 457538 132466 457774
rect 132702 457538 132734 457774
rect 132114 457454 132734 457538
rect 132114 457218 132146 457454
rect 132382 457218 132466 457454
rect 132702 457218 132734 457454
rect 132114 421774 132734 457218
rect 132114 421538 132146 421774
rect 132382 421538 132466 421774
rect 132702 421538 132734 421774
rect 132114 421454 132734 421538
rect 132114 421218 132146 421454
rect 132382 421218 132466 421454
rect 132702 421218 132734 421454
rect 132114 385774 132734 421218
rect 132114 385538 132146 385774
rect 132382 385538 132466 385774
rect 132702 385538 132734 385774
rect 132114 385454 132734 385538
rect 132114 385218 132146 385454
rect 132382 385218 132466 385454
rect 132702 385218 132734 385454
rect 132114 349774 132734 385218
rect 132114 349538 132146 349774
rect 132382 349538 132466 349774
rect 132702 349538 132734 349774
rect 132114 349454 132734 349538
rect 132114 349218 132146 349454
rect 132382 349218 132466 349454
rect 132702 349218 132734 349454
rect 132114 313774 132734 349218
rect 132114 313538 132146 313774
rect 132382 313538 132466 313774
rect 132702 313538 132734 313774
rect 132114 313454 132734 313538
rect 132114 313218 132146 313454
rect 132382 313218 132466 313454
rect 132702 313218 132734 313454
rect 132114 277774 132734 313218
rect 132114 277538 132146 277774
rect 132382 277538 132466 277774
rect 132702 277538 132734 277774
rect 132114 277454 132734 277538
rect 132114 277218 132146 277454
rect 132382 277218 132466 277454
rect 132702 277218 132734 277454
rect 132114 241774 132734 277218
rect 132114 241538 132146 241774
rect 132382 241538 132466 241774
rect 132702 241538 132734 241774
rect 132114 241454 132734 241538
rect 132114 241218 132146 241454
rect 132382 241218 132466 241454
rect 132702 241218 132734 241454
rect 132114 205774 132734 241218
rect 132114 205538 132146 205774
rect 132382 205538 132466 205774
rect 132702 205538 132734 205774
rect 132114 205454 132734 205538
rect 132114 205218 132146 205454
rect 132382 205218 132466 205454
rect 132702 205218 132734 205454
rect 132114 169774 132734 205218
rect 132114 169538 132146 169774
rect 132382 169538 132466 169774
rect 132702 169538 132734 169774
rect 132114 169454 132734 169538
rect 132114 169218 132146 169454
rect 132382 169218 132466 169454
rect 132702 169218 132734 169454
rect 132114 133774 132734 169218
rect 132114 133538 132146 133774
rect 132382 133538 132466 133774
rect 132702 133538 132734 133774
rect 132114 133454 132734 133538
rect 132114 133218 132146 133454
rect 132382 133218 132466 133454
rect 132702 133218 132734 133454
rect 132114 97774 132734 133218
rect 132114 97538 132146 97774
rect 132382 97538 132466 97774
rect 132702 97538 132734 97774
rect 132114 97454 132734 97538
rect 132114 97218 132146 97454
rect 132382 97218 132466 97454
rect 132702 97218 132734 97454
rect 132114 61774 132734 97218
rect 132114 61538 132146 61774
rect 132382 61538 132466 61774
rect 132702 61538 132734 61774
rect 132114 61454 132734 61538
rect 132114 61218 132146 61454
rect 132382 61218 132466 61454
rect 132702 61218 132734 61454
rect 132114 25774 132734 61218
rect 132114 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 132734 25774
rect 132114 25454 132734 25538
rect 132114 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 132734 25454
rect 132114 -6106 132734 25218
rect 132114 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 132734 -6106
rect 132114 -6426 132734 -6342
rect 132114 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 132734 -6426
rect 132114 -7654 132734 -6662
rect 135834 711558 136454 711590
rect 135834 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 136454 711558
rect 135834 711238 136454 711322
rect 135834 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 136454 711238
rect 135834 677494 136454 711002
rect 135834 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 136454 677494
rect 135834 677174 136454 677258
rect 135834 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 136454 677174
rect 135834 641494 136454 676938
rect 135834 641258 135866 641494
rect 136102 641258 136186 641494
rect 136422 641258 136454 641494
rect 135834 641174 136454 641258
rect 135834 640938 135866 641174
rect 136102 640938 136186 641174
rect 136422 640938 136454 641174
rect 135834 605494 136454 640938
rect 135834 605258 135866 605494
rect 136102 605258 136186 605494
rect 136422 605258 136454 605494
rect 135834 605174 136454 605258
rect 135834 604938 135866 605174
rect 136102 604938 136186 605174
rect 136422 604938 136454 605174
rect 135834 569494 136454 604938
rect 135834 569258 135866 569494
rect 136102 569258 136186 569494
rect 136422 569258 136454 569494
rect 135834 569174 136454 569258
rect 135834 568938 135866 569174
rect 136102 568938 136186 569174
rect 136422 568938 136454 569174
rect 135834 533494 136454 568938
rect 135834 533258 135866 533494
rect 136102 533258 136186 533494
rect 136422 533258 136454 533494
rect 135834 533174 136454 533258
rect 135834 532938 135866 533174
rect 136102 532938 136186 533174
rect 136422 532938 136454 533174
rect 135834 497494 136454 532938
rect 135834 497258 135866 497494
rect 136102 497258 136186 497494
rect 136422 497258 136454 497494
rect 135834 497174 136454 497258
rect 135834 496938 135866 497174
rect 136102 496938 136186 497174
rect 136422 496938 136454 497174
rect 135834 461494 136454 496938
rect 135834 461258 135866 461494
rect 136102 461258 136186 461494
rect 136422 461258 136454 461494
rect 135834 461174 136454 461258
rect 135834 460938 135866 461174
rect 136102 460938 136186 461174
rect 136422 460938 136454 461174
rect 135834 425494 136454 460938
rect 135834 425258 135866 425494
rect 136102 425258 136186 425494
rect 136422 425258 136454 425494
rect 135834 425174 136454 425258
rect 135834 424938 135866 425174
rect 136102 424938 136186 425174
rect 136422 424938 136454 425174
rect 135834 389494 136454 424938
rect 135834 389258 135866 389494
rect 136102 389258 136186 389494
rect 136422 389258 136454 389494
rect 135834 389174 136454 389258
rect 135834 388938 135866 389174
rect 136102 388938 136186 389174
rect 136422 388938 136454 389174
rect 135834 353494 136454 388938
rect 135834 353258 135866 353494
rect 136102 353258 136186 353494
rect 136422 353258 136454 353494
rect 135834 353174 136454 353258
rect 135834 352938 135866 353174
rect 136102 352938 136186 353174
rect 136422 352938 136454 353174
rect 135834 317494 136454 352938
rect 135834 317258 135866 317494
rect 136102 317258 136186 317494
rect 136422 317258 136454 317494
rect 135834 317174 136454 317258
rect 135834 316938 135866 317174
rect 136102 316938 136186 317174
rect 136422 316938 136454 317174
rect 135834 281494 136454 316938
rect 135834 281258 135866 281494
rect 136102 281258 136186 281494
rect 136422 281258 136454 281494
rect 135834 281174 136454 281258
rect 135834 280938 135866 281174
rect 136102 280938 136186 281174
rect 136422 280938 136454 281174
rect 135834 245494 136454 280938
rect 135834 245258 135866 245494
rect 136102 245258 136186 245494
rect 136422 245258 136454 245494
rect 135834 245174 136454 245258
rect 135834 244938 135866 245174
rect 136102 244938 136186 245174
rect 136422 244938 136454 245174
rect 135834 209494 136454 244938
rect 135834 209258 135866 209494
rect 136102 209258 136186 209494
rect 136422 209258 136454 209494
rect 135834 209174 136454 209258
rect 135834 208938 135866 209174
rect 136102 208938 136186 209174
rect 136422 208938 136454 209174
rect 135834 173494 136454 208938
rect 135834 173258 135866 173494
rect 136102 173258 136186 173494
rect 136422 173258 136454 173494
rect 135834 173174 136454 173258
rect 135834 172938 135866 173174
rect 136102 172938 136186 173174
rect 136422 172938 136454 173174
rect 135834 137494 136454 172938
rect 135834 137258 135866 137494
rect 136102 137258 136186 137494
rect 136422 137258 136454 137494
rect 135834 137174 136454 137258
rect 135834 136938 135866 137174
rect 136102 136938 136186 137174
rect 136422 136938 136454 137174
rect 135834 101494 136454 136938
rect 135834 101258 135866 101494
rect 136102 101258 136186 101494
rect 136422 101258 136454 101494
rect 135834 101174 136454 101258
rect 135834 100938 135866 101174
rect 136102 100938 136186 101174
rect 136422 100938 136454 101174
rect 135834 65494 136454 100938
rect 135834 65258 135866 65494
rect 136102 65258 136186 65494
rect 136422 65258 136454 65494
rect 135834 65174 136454 65258
rect 135834 64938 135866 65174
rect 136102 64938 136186 65174
rect 136422 64938 136454 65174
rect 135834 29494 136454 64938
rect 135834 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 136454 29494
rect 135834 29174 136454 29258
rect 135834 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 136454 29174
rect 135834 -7066 136454 28938
rect 135834 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 136454 -7066
rect 135834 -7386 136454 -7302
rect 135834 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 136454 -7386
rect 135834 -7654 136454 -7622
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 149514 705798 150134 711590
rect 149514 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 150134 705798
rect 149514 705478 150134 705562
rect 149514 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 150134 705478
rect 149514 691174 150134 705242
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -1306 150134 6618
rect 149514 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 150134 -1306
rect 149514 -1626 150134 -1542
rect 149514 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 150134 -1626
rect 149514 -7654 150134 -1862
rect 153234 706758 153854 711590
rect 153234 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 153854 706758
rect 153234 706438 153854 706522
rect 153234 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 153854 706438
rect 153234 694894 153854 706202
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -2266 153854 10338
rect 153234 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 153854 -2266
rect 153234 -2586 153854 -2502
rect 153234 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 153854 -2586
rect 153234 -7654 153854 -2822
rect 156954 707718 157574 711590
rect 156954 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 157574 707718
rect 156954 707398 157574 707482
rect 156954 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 157574 707398
rect 156954 698614 157574 707162
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 156954 -3226 157574 14058
rect 156954 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 157574 -3226
rect 156954 -3546 157574 -3462
rect 156954 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 157574 -3546
rect 156954 -7654 157574 -3782
rect 160674 708678 161294 711590
rect 160674 708442 160706 708678
rect 160942 708442 161026 708678
rect 161262 708442 161294 708678
rect 160674 708358 161294 708442
rect 160674 708122 160706 708358
rect 160942 708122 161026 708358
rect 161262 708122 161294 708358
rect 160674 666334 161294 708122
rect 160674 666098 160706 666334
rect 160942 666098 161026 666334
rect 161262 666098 161294 666334
rect 160674 666014 161294 666098
rect 160674 665778 160706 666014
rect 160942 665778 161026 666014
rect 161262 665778 161294 666014
rect 160674 630334 161294 665778
rect 160674 630098 160706 630334
rect 160942 630098 161026 630334
rect 161262 630098 161294 630334
rect 160674 630014 161294 630098
rect 160674 629778 160706 630014
rect 160942 629778 161026 630014
rect 161262 629778 161294 630014
rect 160674 594334 161294 629778
rect 160674 594098 160706 594334
rect 160942 594098 161026 594334
rect 161262 594098 161294 594334
rect 160674 594014 161294 594098
rect 160674 593778 160706 594014
rect 160942 593778 161026 594014
rect 161262 593778 161294 594014
rect 160674 558334 161294 593778
rect 160674 558098 160706 558334
rect 160942 558098 161026 558334
rect 161262 558098 161294 558334
rect 160674 558014 161294 558098
rect 160674 557778 160706 558014
rect 160942 557778 161026 558014
rect 161262 557778 161294 558014
rect 160674 522334 161294 557778
rect 160674 522098 160706 522334
rect 160942 522098 161026 522334
rect 161262 522098 161294 522334
rect 160674 522014 161294 522098
rect 160674 521778 160706 522014
rect 160942 521778 161026 522014
rect 161262 521778 161294 522014
rect 160674 486334 161294 521778
rect 160674 486098 160706 486334
rect 160942 486098 161026 486334
rect 161262 486098 161294 486334
rect 160674 486014 161294 486098
rect 160674 485778 160706 486014
rect 160942 485778 161026 486014
rect 161262 485778 161294 486014
rect 160674 450334 161294 485778
rect 160674 450098 160706 450334
rect 160942 450098 161026 450334
rect 161262 450098 161294 450334
rect 160674 450014 161294 450098
rect 160674 449778 160706 450014
rect 160942 449778 161026 450014
rect 161262 449778 161294 450014
rect 160674 414334 161294 449778
rect 160674 414098 160706 414334
rect 160942 414098 161026 414334
rect 161262 414098 161294 414334
rect 160674 414014 161294 414098
rect 160674 413778 160706 414014
rect 160942 413778 161026 414014
rect 161262 413778 161294 414014
rect 160674 378334 161294 413778
rect 160674 378098 160706 378334
rect 160942 378098 161026 378334
rect 161262 378098 161294 378334
rect 160674 378014 161294 378098
rect 160674 377778 160706 378014
rect 160942 377778 161026 378014
rect 161262 377778 161294 378014
rect 160674 342334 161294 377778
rect 160674 342098 160706 342334
rect 160942 342098 161026 342334
rect 161262 342098 161294 342334
rect 160674 342014 161294 342098
rect 160674 341778 160706 342014
rect 160942 341778 161026 342014
rect 161262 341778 161294 342014
rect 160674 306334 161294 341778
rect 160674 306098 160706 306334
rect 160942 306098 161026 306334
rect 161262 306098 161294 306334
rect 160674 306014 161294 306098
rect 160674 305778 160706 306014
rect 160942 305778 161026 306014
rect 161262 305778 161294 306014
rect 160674 270334 161294 305778
rect 160674 270098 160706 270334
rect 160942 270098 161026 270334
rect 161262 270098 161294 270334
rect 160674 270014 161294 270098
rect 160674 269778 160706 270014
rect 160942 269778 161026 270014
rect 161262 269778 161294 270014
rect 160674 234334 161294 269778
rect 160674 234098 160706 234334
rect 160942 234098 161026 234334
rect 161262 234098 161294 234334
rect 160674 234014 161294 234098
rect 160674 233778 160706 234014
rect 160942 233778 161026 234014
rect 161262 233778 161294 234014
rect 160674 198334 161294 233778
rect 160674 198098 160706 198334
rect 160942 198098 161026 198334
rect 161262 198098 161294 198334
rect 160674 198014 161294 198098
rect 160674 197778 160706 198014
rect 160942 197778 161026 198014
rect 161262 197778 161294 198014
rect 160674 162334 161294 197778
rect 160674 162098 160706 162334
rect 160942 162098 161026 162334
rect 161262 162098 161294 162334
rect 160674 162014 161294 162098
rect 160674 161778 160706 162014
rect 160942 161778 161026 162014
rect 161262 161778 161294 162014
rect 160674 126334 161294 161778
rect 160674 126098 160706 126334
rect 160942 126098 161026 126334
rect 161262 126098 161294 126334
rect 160674 126014 161294 126098
rect 160674 125778 160706 126014
rect 160942 125778 161026 126014
rect 161262 125778 161294 126014
rect 160674 90334 161294 125778
rect 160674 90098 160706 90334
rect 160942 90098 161026 90334
rect 161262 90098 161294 90334
rect 160674 90014 161294 90098
rect 160674 89778 160706 90014
rect 160942 89778 161026 90014
rect 161262 89778 161294 90014
rect 160674 54334 161294 89778
rect 160674 54098 160706 54334
rect 160942 54098 161026 54334
rect 161262 54098 161294 54334
rect 160674 54014 161294 54098
rect 160674 53778 160706 54014
rect 160942 53778 161026 54014
rect 161262 53778 161294 54014
rect 160674 18334 161294 53778
rect 160674 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 161294 18334
rect 160674 18014 161294 18098
rect 160674 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 161294 18014
rect 160674 -4186 161294 17778
rect 160674 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 161294 -4186
rect 160674 -4506 161294 -4422
rect 160674 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 161294 -4506
rect 160674 -7654 161294 -4742
rect 164394 709638 165014 711590
rect 164394 709402 164426 709638
rect 164662 709402 164746 709638
rect 164982 709402 165014 709638
rect 164394 709318 165014 709402
rect 164394 709082 164426 709318
rect 164662 709082 164746 709318
rect 164982 709082 165014 709318
rect 164394 670054 165014 709082
rect 164394 669818 164426 670054
rect 164662 669818 164746 670054
rect 164982 669818 165014 670054
rect 164394 669734 165014 669818
rect 164394 669498 164426 669734
rect 164662 669498 164746 669734
rect 164982 669498 165014 669734
rect 164394 634054 165014 669498
rect 164394 633818 164426 634054
rect 164662 633818 164746 634054
rect 164982 633818 165014 634054
rect 164394 633734 165014 633818
rect 164394 633498 164426 633734
rect 164662 633498 164746 633734
rect 164982 633498 165014 633734
rect 164394 598054 165014 633498
rect 164394 597818 164426 598054
rect 164662 597818 164746 598054
rect 164982 597818 165014 598054
rect 164394 597734 165014 597818
rect 164394 597498 164426 597734
rect 164662 597498 164746 597734
rect 164982 597498 165014 597734
rect 164394 562054 165014 597498
rect 164394 561818 164426 562054
rect 164662 561818 164746 562054
rect 164982 561818 165014 562054
rect 164394 561734 165014 561818
rect 164394 561498 164426 561734
rect 164662 561498 164746 561734
rect 164982 561498 165014 561734
rect 164394 526054 165014 561498
rect 164394 525818 164426 526054
rect 164662 525818 164746 526054
rect 164982 525818 165014 526054
rect 164394 525734 165014 525818
rect 164394 525498 164426 525734
rect 164662 525498 164746 525734
rect 164982 525498 165014 525734
rect 164394 490054 165014 525498
rect 164394 489818 164426 490054
rect 164662 489818 164746 490054
rect 164982 489818 165014 490054
rect 164394 489734 165014 489818
rect 164394 489498 164426 489734
rect 164662 489498 164746 489734
rect 164982 489498 165014 489734
rect 164394 454054 165014 489498
rect 164394 453818 164426 454054
rect 164662 453818 164746 454054
rect 164982 453818 165014 454054
rect 164394 453734 165014 453818
rect 164394 453498 164426 453734
rect 164662 453498 164746 453734
rect 164982 453498 165014 453734
rect 164394 418054 165014 453498
rect 164394 417818 164426 418054
rect 164662 417818 164746 418054
rect 164982 417818 165014 418054
rect 164394 417734 165014 417818
rect 164394 417498 164426 417734
rect 164662 417498 164746 417734
rect 164982 417498 165014 417734
rect 164394 382054 165014 417498
rect 164394 381818 164426 382054
rect 164662 381818 164746 382054
rect 164982 381818 165014 382054
rect 164394 381734 165014 381818
rect 164394 381498 164426 381734
rect 164662 381498 164746 381734
rect 164982 381498 165014 381734
rect 164394 346054 165014 381498
rect 164394 345818 164426 346054
rect 164662 345818 164746 346054
rect 164982 345818 165014 346054
rect 164394 345734 165014 345818
rect 164394 345498 164426 345734
rect 164662 345498 164746 345734
rect 164982 345498 165014 345734
rect 164394 310054 165014 345498
rect 164394 309818 164426 310054
rect 164662 309818 164746 310054
rect 164982 309818 165014 310054
rect 164394 309734 165014 309818
rect 164394 309498 164426 309734
rect 164662 309498 164746 309734
rect 164982 309498 165014 309734
rect 164394 274054 165014 309498
rect 164394 273818 164426 274054
rect 164662 273818 164746 274054
rect 164982 273818 165014 274054
rect 164394 273734 165014 273818
rect 164394 273498 164426 273734
rect 164662 273498 164746 273734
rect 164982 273498 165014 273734
rect 164394 238054 165014 273498
rect 164394 237818 164426 238054
rect 164662 237818 164746 238054
rect 164982 237818 165014 238054
rect 164394 237734 165014 237818
rect 164394 237498 164426 237734
rect 164662 237498 164746 237734
rect 164982 237498 165014 237734
rect 164394 202054 165014 237498
rect 168114 710598 168734 711590
rect 168114 710362 168146 710598
rect 168382 710362 168466 710598
rect 168702 710362 168734 710598
rect 168114 710278 168734 710362
rect 168114 710042 168146 710278
rect 168382 710042 168466 710278
rect 168702 710042 168734 710278
rect 168114 673774 168734 710042
rect 168114 673538 168146 673774
rect 168382 673538 168466 673774
rect 168702 673538 168734 673774
rect 168114 673454 168734 673538
rect 168114 673218 168146 673454
rect 168382 673218 168466 673454
rect 168702 673218 168734 673454
rect 168114 637774 168734 673218
rect 168114 637538 168146 637774
rect 168382 637538 168466 637774
rect 168702 637538 168734 637774
rect 168114 637454 168734 637538
rect 168114 637218 168146 637454
rect 168382 637218 168466 637454
rect 168702 637218 168734 637454
rect 168114 601774 168734 637218
rect 168114 601538 168146 601774
rect 168382 601538 168466 601774
rect 168702 601538 168734 601774
rect 168114 601454 168734 601538
rect 168114 601218 168146 601454
rect 168382 601218 168466 601454
rect 168702 601218 168734 601454
rect 168114 565774 168734 601218
rect 168114 565538 168146 565774
rect 168382 565538 168466 565774
rect 168702 565538 168734 565774
rect 168114 565454 168734 565538
rect 168114 565218 168146 565454
rect 168382 565218 168466 565454
rect 168702 565218 168734 565454
rect 168114 529774 168734 565218
rect 168114 529538 168146 529774
rect 168382 529538 168466 529774
rect 168702 529538 168734 529774
rect 168114 529454 168734 529538
rect 168114 529218 168146 529454
rect 168382 529218 168466 529454
rect 168702 529218 168734 529454
rect 168114 493774 168734 529218
rect 168114 493538 168146 493774
rect 168382 493538 168466 493774
rect 168702 493538 168734 493774
rect 168114 493454 168734 493538
rect 168114 493218 168146 493454
rect 168382 493218 168466 493454
rect 168702 493218 168734 493454
rect 168114 457774 168734 493218
rect 168114 457538 168146 457774
rect 168382 457538 168466 457774
rect 168702 457538 168734 457774
rect 168114 457454 168734 457538
rect 168114 457218 168146 457454
rect 168382 457218 168466 457454
rect 168702 457218 168734 457454
rect 168114 421774 168734 457218
rect 168114 421538 168146 421774
rect 168382 421538 168466 421774
rect 168702 421538 168734 421774
rect 168114 421454 168734 421538
rect 168114 421218 168146 421454
rect 168382 421218 168466 421454
rect 168702 421218 168734 421454
rect 168114 385774 168734 421218
rect 168114 385538 168146 385774
rect 168382 385538 168466 385774
rect 168702 385538 168734 385774
rect 168114 385454 168734 385538
rect 168114 385218 168146 385454
rect 168382 385218 168466 385454
rect 168702 385218 168734 385454
rect 168114 349774 168734 385218
rect 168114 349538 168146 349774
rect 168382 349538 168466 349774
rect 168702 349538 168734 349774
rect 168114 349454 168734 349538
rect 168114 349218 168146 349454
rect 168382 349218 168466 349454
rect 168702 349218 168734 349454
rect 168114 313774 168734 349218
rect 168114 313538 168146 313774
rect 168382 313538 168466 313774
rect 168702 313538 168734 313774
rect 168114 313454 168734 313538
rect 168114 313218 168146 313454
rect 168382 313218 168466 313454
rect 168702 313218 168734 313454
rect 168114 277774 168734 313218
rect 168114 277538 168146 277774
rect 168382 277538 168466 277774
rect 168702 277538 168734 277774
rect 168114 277454 168734 277538
rect 168114 277218 168146 277454
rect 168382 277218 168466 277454
rect 168702 277218 168734 277454
rect 168114 241774 168734 277218
rect 168114 241538 168146 241774
rect 168382 241538 168466 241774
rect 168702 241538 168734 241774
rect 168114 241454 168734 241538
rect 168114 241218 168146 241454
rect 168382 241218 168466 241454
rect 168702 241218 168734 241454
rect 167499 217700 167565 217701
rect 167499 217636 167500 217700
rect 167564 217636 167565 217700
rect 167499 217635 167565 217636
rect 167315 204780 167381 204781
rect 167315 204716 167316 204780
rect 167380 204716 167381 204780
rect 167315 204715 167381 204716
rect 164394 201818 164426 202054
rect 164662 201818 164746 202054
rect 164982 201818 165014 202054
rect 164394 201734 165014 201818
rect 164394 201498 164426 201734
rect 164662 201498 164746 201734
rect 164982 201498 165014 201734
rect 164394 166054 165014 201498
rect 164394 165818 164426 166054
rect 164662 165818 164746 166054
rect 164982 165818 165014 166054
rect 164394 165734 165014 165818
rect 164394 165498 164426 165734
rect 164662 165498 164746 165734
rect 164982 165498 165014 165734
rect 164394 130054 165014 165498
rect 164394 129818 164426 130054
rect 164662 129818 164746 130054
rect 164982 129818 165014 130054
rect 164394 129734 165014 129818
rect 164394 129498 164426 129734
rect 164662 129498 164746 129734
rect 164982 129498 165014 129734
rect 164394 94054 165014 129498
rect 166027 119372 166093 119373
rect 166027 119308 166028 119372
rect 166092 119308 166093 119372
rect 166027 119307 166093 119308
rect 166030 118013 166090 119307
rect 166947 118828 167013 118829
rect 166947 118764 166948 118828
rect 167012 118764 167013 118828
rect 166947 118763 167013 118764
rect 166027 118012 166093 118013
rect 166027 117948 166028 118012
rect 166092 117948 166093 118012
rect 166027 117947 166093 117948
rect 166950 116517 167010 118763
rect 166947 116516 167013 116517
rect 166947 116452 166948 116516
rect 167012 116452 167013 116516
rect 166947 116451 167013 116452
rect 167318 111893 167378 204715
rect 167502 112301 167562 217635
rect 168114 205774 168734 241218
rect 171834 711558 172454 711590
rect 171834 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 172454 711558
rect 171834 711238 172454 711322
rect 171834 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 172454 711238
rect 171834 677494 172454 711002
rect 171834 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 172454 677494
rect 171834 677174 172454 677258
rect 171834 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 172454 677174
rect 171834 641494 172454 676938
rect 171834 641258 171866 641494
rect 172102 641258 172186 641494
rect 172422 641258 172454 641494
rect 171834 641174 172454 641258
rect 171834 640938 171866 641174
rect 172102 640938 172186 641174
rect 172422 640938 172454 641174
rect 171834 605494 172454 640938
rect 171834 605258 171866 605494
rect 172102 605258 172186 605494
rect 172422 605258 172454 605494
rect 171834 605174 172454 605258
rect 171834 604938 171866 605174
rect 172102 604938 172186 605174
rect 172422 604938 172454 605174
rect 171834 569494 172454 604938
rect 171834 569258 171866 569494
rect 172102 569258 172186 569494
rect 172422 569258 172454 569494
rect 171834 569174 172454 569258
rect 171834 568938 171866 569174
rect 172102 568938 172186 569174
rect 172422 568938 172454 569174
rect 171834 533494 172454 568938
rect 171834 533258 171866 533494
rect 172102 533258 172186 533494
rect 172422 533258 172454 533494
rect 171834 533174 172454 533258
rect 171834 532938 171866 533174
rect 172102 532938 172186 533174
rect 172422 532938 172454 533174
rect 171834 497494 172454 532938
rect 171834 497258 171866 497494
rect 172102 497258 172186 497494
rect 172422 497258 172454 497494
rect 171834 497174 172454 497258
rect 171834 496938 171866 497174
rect 172102 496938 172186 497174
rect 172422 496938 172454 497174
rect 171834 461494 172454 496938
rect 171834 461258 171866 461494
rect 172102 461258 172186 461494
rect 172422 461258 172454 461494
rect 171834 461174 172454 461258
rect 171834 460938 171866 461174
rect 172102 460938 172186 461174
rect 172422 460938 172454 461174
rect 171834 425494 172454 460938
rect 171834 425258 171866 425494
rect 172102 425258 172186 425494
rect 172422 425258 172454 425494
rect 171834 425174 172454 425258
rect 171834 424938 171866 425174
rect 172102 424938 172186 425174
rect 172422 424938 172454 425174
rect 171834 389494 172454 424938
rect 171834 389258 171866 389494
rect 172102 389258 172186 389494
rect 172422 389258 172454 389494
rect 171834 389174 172454 389258
rect 171834 388938 171866 389174
rect 172102 388938 172186 389174
rect 172422 388938 172454 389174
rect 171834 353494 172454 388938
rect 171834 353258 171866 353494
rect 172102 353258 172186 353494
rect 172422 353258 172454 353494
rect 171834 353174 172454 353258
rect 171834 352938 171866 353174
rect 172102 352938 172186 353174
rect 172422 352938 172454 353174
rect 171834 317494 172454 352938
rect 171834 317258 171866 317494
rect 172102 317258 172186 317494
rect 172422 317258 172454 317494
rect 171834 317174 172454 317258
rect 171834 316938 171866 317174
rect 172102 316938 172186 317174
rect 172422 316938 172454 317174
rect 171834 281494 172454 316938
rect 171834 281258 171866 281494
rect 172102 281258 172186 281494
rect 172422 281258 172454 281494
rect 171834 281174 172454 281258
rect 171834 280938 171866 281174
rect 172102 280938 172186 281174
rect 172422 280938 172454 281174
rect 171834 245494 172454 280938
rect 171834 245258 171866 245494
rect 172102 245258 172186 245494
rect 172422 245258 172454 245494
rect 171834 245174 172454 245258
rect 171834 244938 171866 245174
rect 172102 244938 172186 245174
rect 172422 244938 172454 245174
rect 169523 233884 169589 233885
rect 169523 233820 169524 233884
rect 169588 233820 169589 233884
rect 169523 233819 169589 233820
rect 168114 205538 168146 205774
rect 168382 205538 168466 205774
rect 168702 205538 168734 205774
rect 168114 205454 168734 205538
rect 168114 205218 168146 205454
rect 168382 205218 168466 205454
rect 168702 205218 168734 205454
rect 167683 195260 167749 195261
rect 167683 195196 167684 195260
rect 167748 195196 167749 195260
rect 167683 195195 167749 195196
rect 167499 112300 167565 112301
rect 167499 112236 167500 112300
rect 167564 112236 167565 112300
rect 167499 112235 167565 112236
rect 167315 111892 167381 111893
rect 167315 111828 167316 111892
rect 167380 111828 167381 111892
rect 167315 111827 167381 111828
rect 167502 101285 167562 112235
rect 167499 101284 167565 101285
rect 167499 101220 167500 101284
rect 167564 101220 167565 101284
rect 167499 101219 167565 101220
rect 167499 96524 167565 96525
rect 167499 96460 167500 96524
rect 167564 96460 167565 96524
rect 167499 96459 167565 96460
rect 167315 95844 167381 95845
rect 167315 95780 167316 95844
rect 167380 95780 167381 95844
rect 167315 95779 167381 95780
rect 164394 93818 164426 94054
rect 164662 93818 164746 94054
rect 164982 93818 165014 94054
rect 164394 93734 165014 93818
rect 164394 93498 164426 93734
rect 164662 93498 164746 93734
rect 164982 93498 165014 93734
rect 164394 58054 165014 93498
rect 167318 69733 167378 95779
rect 167315 69732 167381 69733
rect 167315 69668 167316 69732
rect 167380 69668 167381 69732
rect 167315 69667 167381 69668
rect 164394 57818 164426 58054
rect 164662 57818 164746 58054
rect 164982 57818 165014 58054
rect 164394 57734 165014 57818
rect 164394 57498 164426 57734
rect 164662 57498 164746 57734
rect 164982 57498 165014 57734
rect 164394 22054 165014 57498
rect 167502 54501 167562 96459
rect 167686 87549 167746 195195
rect 167867 193220 167933 193221
rect 167867 193156 167868 193220
rect 167932 193156 167933 193220
rect 167867 193155 167933 193156
rect 167683 87548 167749 87549
rect 167683 87484 167684 87548
rect 167748 87484 167749 87548
rect 167683 87483 167749 87484
rect 167870 85101 167930 193155
rect 168114 169774 168734 205218
rect 169526 175541 169586 233819
rect 169707 230620 169773 230621
rect 169707 230556 169708 230620
rect 169772 230556 169773 230620
rect 169707 230555 169773 230556
rect 169523 175540 169589 175541
rect 169523 175476 169524 175540
rect 169588 175476 169589 175540
rect 169523 175475 169589 175476
rect 168114 169538 168146 169774
rect 168382 169538 168466 169774
rect 168702 169538 168734 169774
rect 168114 169454 168734 169538
rect 168114 169218 168146 169454
rect 168382 169218 168466 169454
rect 168702 169218 168734 169454
rect 168114 133774 168734 169218
rect 168114 133538 168146 133774
rect 168382 133538 168466 133774
rect 168702 133538 168734 133774
rect 168114 133454 168734 133538
rect 168114 133218 168146 133454
rect 168382 133218 168466 133454
rect 168702 133218 168734 133454
rect 168114 97774 168734 133218
rect 169710 132510 169770 230555
rect 171834 209494 172454 244938
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 174208 219454 174528 219486
rect 174208 219218 174250 219454
rect 174486 219218 174528 219454
rect 174208 219134 174528 219218
rect 174208 218898 174250 219134
rect 174486 218898 174528 219134
rect 174208 218866 174528 218898
rect 181794 219454 182414 254898
rect 185514 705798 186134 711590
rect 185514 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 186134 705798
rect 185514 705478 186134 705562
rect 185514 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 186134 705478
rect 185514 691174 186134 705242
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 225473 186134 258618
rect 189234 706758 189854 711590
rect 189234 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 189854 706758
rect 189234 706438 189854 706522
rect 189234 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 189854 706438
rect 189234 694894 189854 706202
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 229772 189854 262338
rect 192954 707718 193574 711590
rect 192954 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 193574 707718
rect 192954 707398 193574 707482
rect 192954 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 193574 707398
rect 192954 698614 193574 707162
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 225473 193574 230058
rect 196674 708678 197294 711590
rect 196674 708442 196706 708678
rect 196942 708442 197026 708678
rect 197262 708442 197294 708678
rect 196674 708358 197294 708442
rect 196674 708122 196706 708358
rect 196942 708122 197026 708358
rect 197262 708122 197294 708358
rect 196674 666334 197294 708122
rect 196674 666098 196706 666334
rect 196942 666098 197026 666334
rect 197262 666098 197294 666334
rect 196674 666014 197294 666098
rect 196674 665778 196706 666014
rect 196942 665778 197026 666014
rect 197262 665778 197294 666014
rect 196674 630334 197294 665778
rect 196674 630098 196706 630334
rect 196942 630098 197026 630334
rect 197262 630098 197294 630334
rect 196674 630014 197294 630098
rect 196674 629778 196706 630014
rect 196942 629778 197026 630014
rect 197262 629778 197294 630014
rect 196674 594334 197294 629778
rect 196674 594098 196706 594334
rect 196942 594098 197026 594334
rect 197262 594098 197294 594334
rect 196674 594014 197294 594098
rect 196674 593778 196706 594014
rect 196942 593778 197026 594014
rect 197262 593778 197294 594014
rect 196674 558334 197294 593778
rect 196674 558098 196706 558334
rect 196942 558098 197026 558334
rect 197262 558098 197294 558334
rect 196674 558014 197294 558098
rect 196674 557778 196706 558014
rect 196942 557778 197026 558014
rect 197262 557778 197294 558014
rect 196674 522334 197294 557778
rect 196674 522098 196706 522334
rect 196942 522098 197026 522334
rect 197262 522098 197294 522334
rect 196674 522014 197294 522098
rect 196674 521778 196706 522014
rect 196942 521778 197026 522014
rect 197262 521778 197294 522014
rect 196674 486334 197294 521778
rect 196674 486098 196706 486334
rect 196942 486098 197026 486334
rect 197262 486098 197294 486334
rect 196674 486014 197294 486098
rect 196674 485778 196706 486014
rect 196942 485778 197026 486014
rect 197262 485778 197294 486014
rect 196674 450334 197294 485778
rect 196674 450098 196706 450334
rect 196942 450098 197026 450334
rect 197262 450098 197294 450334
rect 196674 450014 197294 450098
rect 196674 449778 196706 450014
rect 196942 449778 197026 450014
rect 197262 449778 197294 450014
rect 196674 414334 197294 449778
rect 196674 414098 196706 414334
rect 196942 414098 197026 414334
rect 197262 414098 197294 414334
rect 196674 414014 197294 414098
rect 196674 413778 196706 414014
rect 196942 413778 197026 414014
rect 197262 413778 197294 414014
rect 196674 378334 197294 413778
rect 196674 378098 196706 378334
rect 196942 378098 197026 378334
rect 197262 378098 197294 378334
rect 196674 378014 197294 378098
rect 196674 377778 196706 378014
rect 196942 377778 197026 378014
rect 197262 377778 197294 378014
rect 196674 342334 197294 377778
rect 196674 342098 196706 342334
rect 196942 342098 197026 342334
rect 197262 342098 197294 342334
rect 196674 342014 197294 342098
rect 196674 341778 196706 342014
rect 196942 341778 197026 342014
rect 197262 341778 197294 342014
rect 196674 306334 197294 341778
rect 196674 306098 196706 306334
rect 196942 306098 197026 306334
rect 197262 306098 197294 306334
rect 196674 306014 197294 306098
rect 196674 305778 196706 306014
rect 196942 305778 197026 306014
rect 197262 305778 197294 306014
rect 196674 270334 197294 305778
rect 196674 270098 196706 270334
rect 196942 270098 197026 270334
rect 197262 270098 197294 270334
rect 196674 270014 197294 270098
rect 196674 269778 196706 270014
rect 196942 269778 197026 270014
rect 197262 269778 197294 270014
rect 196674 234334 197294 269778
rect 196674 234098 196706 234334
rect 196942 234098 197026 234334
rect 197262 234098 197294 234334
rect 196674 234014 197294 234098
rect 196674 233778 196706 234014
rect 196942 233778 197026 234014
rect 197262 233778 197294 234014
rect 196674 225473 197294 233778
rect 200394 709638 201014 711590
rect 200394 709402 200426 709638
rect 200662 709402 200746 709638
rect 200982 709402 201014 709638
rect 200394 709318 201014 709402
rect 200394 709082 200426 709318
rect 200662 709082 200746 709318
rect 200982 709082 201014 709318
rect 200394 670054 201014 709082
rect 200394 669818 200426 670054
rect 200662 669818 200746 670054
rect 200982 669818 201014 670054
rect 200394 669734 201014 669818
rect 200394 669498 200426 669734
rect 200662 669498 200746 669734
rect 200982 669498 201014 669734
rect 200394 634054 201014 669498
rect 200394 633818 200426 634054
rect 200662 633818 200746 634054
rect 200982 633818 201014 634054
rect 200394 633734 201014 633818
rect 200394 633498 200426 633734
rect 200662 633498 200746 633734
rect 200982 633498 201014 633734
rect 200394 598054 201014 633498
rect 200394 597818 200426 598054
rect 200662 597818 200746 598054
rect 200982 597818 201014 598054
rect 200394 597734 201014 597818
rect 200394 597498 200426 597734
rect 200662 597498 200746 597734
rect 200982 597498 201014 597734
rect 200394 562054 201014 597498
rect 200394 561818 200426 562054
rect 200662 561818 200746 562054
rect 200982 561818 201014 562054
rect 200394 561734 201014 561818
rect 200394 561498 200426 561734
rect 200662 561498 200746 561734
rect 200982 561498 201014 561734
rect 200394 526054 201014 561498
rect 200394 525818 200426 526054
rect 200662 525818 200746 526054
rect 200982 525818 201014 526054
rect 200394 525734 201014 525818
rect 200394 525498 200426 525734
rect 200662 525498 200746 525734
rect 200982 525498 201014 525734
rect 200394 490054 201014 525498
rect 200394 489818 200426 490054
rect 200662 489818 200746 490054
rect 200982 489818 201014 490054
rect 200394 489734 201014 489818
rect 200394 489498 200426 489734
rect 200662 489498 200746 489734
rect 200982 489498 201014 489734
rect 200394 454054 201014 489498
rect 200394 453818 200426 454054
rect 200662 453818 200746 454054
rect 200982 453818 201014 454054
rect 200394 453734 201014 453818
rect 200394 453498 200426 453734
rect 200662 453498 200746 453734
rect 200982 453498 201014 453734
rect 200394 418054 201014 453498
rect 200394 417818 200426 418054
rect 200662 417818 200746 418054
rect 200982 417818 201014 418054
rect 200394 417734 201014 417818
rect 200394 417498 200426 417734
rect 200662 417498 200746 417734
rect 200982 417498 201014 417734
rect 200394 382054 201014 417498
rect 200394 381818 200426 382054
rect 200662 381818 200746 382054
rect 200982 381818 201014 382054
rect 200394 381734 201014 381818
rect 200394 381498 200426 381734
rect 200662 381498 200746 381734
rect 200982 381498 201014 381734
rect 200394 346054 201014 381498
rect 200394 345818 200426 346054
rect 200662 345818 200746 346054
rect 200982 345818 201014 346054
rect 200394 345734 201014 345818
rect 200394 345498 200426 345734
rect 200662 345498 200746 345734
rect 200982 345498 201014 345734
rect 200394 310054 201014 345498
rect 200394 309818 200426 310054
rect 200662 309818 200746 310054
rect 200982 309818 201014 310054
rect 200394 309734 201014 309818
rect 200394 309498 200426 309734
rect 200662 309498 200746 309734
rect 200982 309498 201014 309734
rect 200394 274054 201014 309498
rect 200394 273818 200426 274054
rect 200662 273818 200746 274054
rect 200982 273818 201014 274054
rect 200394 273734 201014 273818
rect 200394 273498 200426 273734
rect 200662 273498 200746 273734
rect 200982 273498 201014 273734
rect 200394 238054 201014 273498
rect 200394 237818 200426 238054
rect 200662 237818 200746 238054
rect 200982 237818 201014 238054
rect 200394 237734 201014 237818
rect 200394 237498 200426 237734
rect 200662 237498 200746 237734
rect 200982 237498 201014 237734
rect 200394 225473 201014 237498
rect 204114 710598 204734 711590
rect 204114 710362 204146 710598
rect 204382 710362 204466 710598
rect 204702 710362 204734 710598
rect 204114 710278 204734 710362
rect 204114 710042 204146 710278
rect 204382 710042 204466 710278
rect 204702 710042 204734 710278
rect 204114 673774 204734 710042
rect 204114 673538 204146 673774
rect 204382 673538 204466 673774
rect 204702 673538 204734 673774
rect 204114 673454 204734 673538
rect 204114 673218 204146 673454
rect 204382 673218 204466 673454
rect 204702 673218 204734 673454
rect 204114 637774 204734 673218
rect 204114 637538 204146 637774
rect 204382 637538 204466 637774
rect 204702 637538 204734 637774
rect 204114 637454 204734 637538
rect 204114 637218 204146 637454
rect 204382 637218 204466 637454
rect 204702 637218 204734 637454
rect 204114 601774 204734 637218
rect 204114 601538 204146 601774
rect 204382 601538 204466 601774
rect 204702 601538 204734 601774
rect 204114 601454 204734 601538
rect 204114 601218 204146 601454
rect 204382 601218 204466 601454
rect 204702 601218 204734 601454
rect 204114 565774 204734 601218
rect 204114 565538 204146 565774
rect 204382 565538 204466 565774
rect 204702 565538 204734 565774
rect 204114 565454 204734 565538
rect 204114 565218 204146 565454
rect 204382 565218 204466 565454
rect 204702 565218 204734 565454
rect 204114 529774 204734 565218
rect 204114 529538 204146 529774
rect 204382 529538 204466 529774
rect 204702 529538 204734 529774
rect 204114 529454 204734 529538
rect 204114 529218 204146 529454
rect 204382 529218 204466 529454
rect 204702 529218 204734 529454
rect 204114 493774 204734 529218
rect 204114 493538 204146 493774
rect 204382 493538 204466 493774
rect 204702 493538 204734 493774
rect 204114 493454 204734 493538
rect 204114 493218 204146 493454
rect 204382 493218 204466 493454
rect 204702 493218 204734 493454
rect 204114 457774 204734 493218
rect 204114 457538 204146 457774
rect 204382 457538 204466 457774
rect 204702 457538 204734 457774
rect 204114 457454 204734 457538
rect 204114 457218 204146 457454
rect 204382 457218 204466 457454
rect 204702 457218 204734 457454
rect 204114 421774 204734 457218
rect 204114 421538 204146 421774
rect 204382 421538 204466 421774
rect 204702 421538 204734 421774
rect 204114 421454 204734 421538
rect 204114 421218 204146 421454
rect 204382 421218 204466 421454
rect 204702 421218 204734 421454
rect 204114 385774 204734 421218
rect 204114 385538 204146 385774
rect 204382 385538 204466 385774
rect 204702 385538 204734 385774
rect 204114 385454 204734 385538
rect 204114 385218 204146 385454
rect 204382 385218 204466 385454
rect 204702 385218 204734 385454
rect 204114 349774 204734 385218
rect 204114 349538 204146 349774
rect 204382 349538 204466 349774
rect 204702 349538 204734 349774
rect 204114 349454 204734 349538
rect 204114 349218 204146 349454
rect 204382 349218 204466 349454
rect 204702 349218 204734 349454
rect 204114 313774 204734 349218
rect 204114 313538 204146 313774
rect 204382 313538 204466 313774
rect 204702 313538 204734 313774
rect 204114 313454 204734 313538
rect 204114 313218 204146 313454
rect 204382 313218 204466 313454
rect 204702 313218 204734 313454
rect 204114 277774 204734 313218
rect 204114 277538 204146 277774
rect 204382 277538 204466 277774
rect 204702 277538 204734 277774
rect 204114 277454 204734 277538
rect 204114 277218 204146 277454
rect 204382 277218 204466 277454
rect 204702 277218 204734 277454
rect 204114 241774 204734 277218
rect 204114 241538 204146 241774
rect 204382 241538 204466 241774
rect 204702 241538 204734 241774
rect 204114 241454 204734 241538
rect 204114 241218 204146 241454
rect 204382 241218 204466 241454
rect 204702 241218 204734 241454
rect 204114 225473 204734 241218
rect 207834 711558 208454 711590
rect 207834 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 208454 711558
rect 207834 711238 208454 711322
rect 207834 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 208454 711238
rect 207834 677494 208454 711002
rect 207834 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 208454 677494
rect 207834 677174 208454 677258
rect 207834 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 208454 677174
rect 207834 641494 208454 676938
rect 207834 641258 207866 641494
rect 208102 641258 208186 641494
rect 208422 641258 208454 641494
rect 207834 641174 208454 641258
rect 207834 640938 207866 641174
rect 208102 640938 208186 641174
rect 208422 640938 208454 641174
rect 207834 605494 208454 640938
rect 207834 605258 207866 605494
rect 208102 605258 208186 605494
rect 208422 605258 208454 605494
rect 207834 605174 208454 605258
rect 207834 604938 207866 605174
rect 208102 604938 208186 605174
rect 208422 604938 208454 605174
rect 207834 569494 208454 604938
rect 207834 569258 207866 569494
rect 208102 569258 208186 569494
rect 208422 569258 208454 569494
rect 207834 569174 208454 569258
rect 207834 568938 207866 569174
rect 208102 568938 208186 569174
rect 208422 568938 208454 569174
rect 207834 533494 208454 568938
rect 207834 533258 207866 533494
rect 208102 533258 208186 533494
rect 208422 533258 208454 533494
rect 207834 533174 208454 533258
rect 207834 532938 207866 533174
rect 208102 532938 208186 533174
rect 208422 532938 208454 533174
rect 207834 497494 208454 532938
rect 207834 497258 207866 497494
rect 208102 497258 208186 497494
rect 208422 497258 208454 497494
rect 207834 497174 208454 497258
rect 207834 496938 207866 497174
rect 208102 496938 208186 497174
rect 208422 496938 208454 497174
rect 207834 461494 208454 496938
rect 207834 461258 207866 461494
rect 208102 461258 208186 461494
rect 208422 461258 208454 461494
rect 207834 461174 208454 461258
rect 207834 460938 207866 461174
rect 208102 460938 208186 461174
rect 208422 460938 208454 461174
rect 207834 425494 208454 460938
rect 207834 425258 207866 425494
rect 208102 425258 208186 425494
rect 208422 425258 208454 425494
rect 207834 425174 208454 425258
rect 207834 424938 207866 425174
rect 208102 424938 208186 425174
rect 208422 424938 208454 425174
rect 207834 389494 208454 424938
rect 207834 389258 207866 389494
rect 208102 389258 208186 389494
rect 208422 389258 208454 389494
rect 207834 389174 208454 389258
rect 207834 388938 207866 389174
rect 208102 388938 208186 389174
rect 208422 388938 208454 389174
rect 207834 353494 208454 388938
rect 207834 353258 207866 353494
rect 208102 353258 208186 353494
rect 208422 353258 208454 353494
rect 207834 353174 208454 353258
rect 207834 352938 207866 353174
rect 208102 352938 208186 353174
rect 208422 352938 208454 353174
rect 207834 317494 208454 352938
rect 207834 317258 207866 317494
rect 208102 317258 208186 317494
rect 208422 317258 208454 317494
rect 207834 317174 208454 317258
rect 207834 316938 207866 317174
rect 208102 316938 208186 317174
rect 208422 316938 208454 317174
rect 207834 281494 208454 316938
rect 207834 281258 207866 281494
rect 208102 281258 208186 281494
rect 208422 281258 208454 281494
rect 207834 281174 208454 281258
rect 207834 280938 207866 281174
rect 208102 280938 208186 281174
rect 208422 280938 208454 281174
rect 207834 245494 208454 280938
rect 207834 245258 207866 245494
rect 208102 245258 208186 245494
rect 208422 245258 208454 245494
rect 207834 245174 208454 245258
rect 207834 244938 207866 245174
rect 208102 244938 208186 245174
rect 208422 244938 208454 245174
rect 207834 225473 208454 244938
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 225473 218414 254898
rect 221514 705798 222134 711590
rect 221514 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 222134 705798
rect 221514 705478 222134 705562
rect 221514 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 222134 705478
rect 221514 691174 222134 705242
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 189568 223174 189888 223206
rect 189568 222938 189610 223174
rect 189846 222938 189888 223174
rect 189568 222854 189888 222938
rect 189568 222618 189610 222854
rect 189846 222618 189888 222854
rect 189568 222586 189888 222618
rect 220288 223174 220608 223206
rect 220288 222938 220330 223174
rect 220566 222938 220608 223174
rect 220288 222854 220608 222938
rect 220288 222618 220330 222854
rect 220566 222618 220608 222854
rect 220288 222586 220608 222618
rect 221514 223174 222134 258618
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 171834 209258 171866 209494
rect 172102 209258 172186 209494
rect 172422 209258 172454 209494
rect 171834 209174 172454 209258
rect 171834 208938 171866 209174
rect 172102 208938 172186 209174
rect 172422 208938 172454 209174
rect 169891 198388 169957 198389
rect 169891 198324 169892 198388
rect 169956 198324 169957 198388
rect 169891 198323 169957 198324
rect 169894 169557 169954 198323
rect 171834 173494 172454 208938
rect 174208 183454 174528 183486
rect 174208 183218 174250 183454
rect 174486 183218 174528 183454
rect 174208 183134 174528 183218
rect 174208 182898 174250 183134
rect 174486 182898 174528 183134
rect 174208 182866 174528 182898
rect 181794 183454 182414 218898
rect 204928 219454 205248 219486
rect 204928 219218 204970 219454
rect 205206 219218 205248 219454
rect 204928 219134 205248 219218
rect 204928 218898 204970 219134
rect 205206 218898 205248 219134
rect 204928 218866 205248 218898
rect 189568 187174 189888 187206
rect 189568 186938 189610 187174
rect 189846 186938 189888 187174
rect 189568 186854 189888 186938
rect 189568 186618 189610 186854
rect 189846 186618 189888 186854
rect 189568 186586 189888 186618
rect 220288 187174 220608 187206
rect 220288 186938 220330 187174
rect 220566 186938 220608 187174
rect 220288 186854 220608 186938
rect 220288 186618 220330 186854
rect 220566 186618 220608 186854
rect 220288 186586 220608 186618
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 171834 173258 171866 173494
rect 172102 173258 172186 173494
rect 172422 173258 172454 173494
rect 171834 173174 172454 173258
rect 171834 172938 171866 173174
rect 172102 172938 172186 173174
rect 172422 172938 172454 173174
rect 169891 169556 169957 169557
rect 169891 169492 169892 169556
rect 169956 169492 169957 169556
rect 169891 169491 169957 169492
rect 171834 137494 172454 172938
rect 171834 137258 171866 137494
rect 172102 137258 172186 137494
rect 172422 137258 172454 137494
rect 171834 137174 172454 137258
rect 171834 136938 171866 137174
rect 172102 136938 172186 137174
rect 172422 136938 172454 137174
rect 169710 132450 170322 132510
rect 170075 120732 170141 120733
rect 170075 120668 170076 120732
rect 170140 120668 170141 120732
rect 170075 120667 170141 120668
rect 169891 120460 169957 120461
rect 169891 120396 169892 120460
rect 169956 120396 169957 120460
rect 169891 120395 169957 120396
rect 169707 120188 169773 120189
rect 169707 120124 169708 120188
rect 169772 120124 169773 120188
rect 169707 120123 169773 120124
rect 169710 113797 169770 120123
rect 169894 113933 169954 120395
rect 170078 114069 170138 120667
rect 170262 116925 170322 132450
rect 170259 116924 170325 116925
rect 170259 116860 170260 116924
rect 170324 116860 170325 116924
rect 170259 116859 170325 116860
rect 170259 114884 170325 114885
rect 170259 114820 170260 114884
rect 170324 114820 170325 114884
rect 170259 114819 170325 114820
rect 170075 114068 170141 114069
rect 170075 114004 170076 114068
rect 170140 114004 170141 114068
rect 170075 114003 170141 114004
rect 169891 113932 169957 113933
rect 169891 113868 169892 113932
rect 169956 113868 169957 113932
rect 169891 113867 169957 113868
rect 169707 113796 169773 113797
rect 169707 113732 169708 113796
rect 169772 113732 169773 113796
rect 169707 113731 169773 113732
rect 170262 113190 170322 114819
rect 169710 113130 170322 113190
rect 169339 110804 169405 110805
rect 169339 110740 169340 110804
rect 169404 110740 169405 110804
rect 169339 110739 169405 110740
rect 168114 97538 168146 97774
rect 168382 97538 168466 97774
rect 168702 97538 168734 97774
rect 168114 97454 168734 97538
rect 168114 97218 168146 97454
rect 168382 97218 168466 97454
rect 168702 97218 168734 97454
rect 167867 85100 167933 85101
rect 167867 85036 167868 85100
rect 167932 85036 167933 85100
rect 167867 85035 167933 85036
rect 167870 84210 167930 85035
rect 167686 84150 167930 84210
rect 167686 69869 167746 84150
rect 167867 72724 167933 72725
rect 167867 72660 167868 72724
rect 167932 72660 167933 72724
rect 167867 72659 167933 72660
rect 167683 69868 167749 69869
rect 167683 69804 167684 69868
rect 167748 69804 167749 69868
rect 167683 69803 167749 69804
rect 167870 64837 167930 72659
rect 167867 64836 167933 64837
rect 167867 64772 167868 64836
rect 167932 64772 167933 64836
rect 167867 64771 167933 64772
rect 167870 58581 167930 64771
rect 168114 61774 168734 97218
rect 168971 73948 169037 73949
rect 168971 73884 168972 73948
rect 169036 73884 169037 73948
rect 168971 73883 169037 73884
rect 168974 69869 169034 73883
rect 168971 69868 169037 69869
rect 168971 69804 168972 69868
rect 169036 69804 169037 69868
rect 168971 69803 169037 69804
rect 168114 61538 168146 61774
rect 168382 61538 168466 61774
rect 168702 61538 168734 61774
rect 168114 61454 168734 61538
rect 168114 61218 168146 61454
rect 168382 61218 168466 61454
rect 168702 61218 168734 61454
rect 167867 58580 167933 58581
rect 167867 58516 167868 58580
rect 167932 58516 167933 58580
rect 167867 58515 167933 58516
rect 167499 54500 167565 54501
rect 167499 54436 167500 54500
rect 167564 54436 167565 54500
rect 167499 54435 167565 54436
rect 164394 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 165014 22054
rect 164394 21734 165014 21818
rect 164394 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 165014 21734
rect 164394 -5146 165014 21498
rect 164394 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 165014 -5146
rect 164394 -5466 165014 -5382
rect 164394 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 165014 -5466
rect 164394 -7654 165014 -5702
rect 168114 25774 168734 61218
rect 169342 53141 169402 110739
rect 169523 101284 169589 101285
rect 169523 101220 169524 101284
rect 169588 101220 169589 101284
rect 169523 101219 169589 101220
rect 169339 53140 169405 53141
rect 169339 53076 169340 53140
rect 169404 53076 169405 53140
rect 169339 53075 169405 53076
rect 168114 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 168734 25774
rect 168114 25454 168734 25538
rect 168114 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 168734 25454
rect 168114 -6106 168734 25218
rect 169526 19957 169586 101219
rect 169710 43485 169770 113130
rect 169891 108900 169957 108901
rect 169891 108836 169892 108900
rect 169956 108836 169957 108900
rect 169891 108835 169957 108836
rect 169707 43484 169773 43485
rect 169707 43420 169708 43484
rect 169772 43420 169773 43484
rect 169707 43419 169773 43420
rect 169894 40629 169954 108835
rect 171834 101494 172454 136938
rect 181794 147454 182414 182898
rect 204928 183454 205248 183486
rect 204928 183218 204970 183454
rect 205206 183218 205248 183454
rect 204928 183134 205248 183218
rect 204928 182898 204970 183134
rect 205206 182898 205248 183134
rect 204928 182866 205248 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 177890 115174 178210 115206
rect 177890 114938 177932 115174
rect 178168 114938 178210 115174
rect 177890 114854 178210 114938
rect 177890 114618 177932 114854
rect 178168 114618 178210 114854
rect 177890 114586 178210 114618
rect 174417 111454 174737 111486
rect 174417 111218 174459 111454
rect 174695 111218 174737 111454
rect 174417 111134 174737 111218
rect 174417 110898 174459 111134
rect 174695 110898 174737 111134
rect 174417 110866 174737 110898
rect 181363 111454 181683 111486
rect 181363 111218 181405 111454
rect 181641 111218 181683 111454
rect 181363 111134 181683 111218
rect 181363 110898 181405 111134
rect 181641 110898 181683 111134
rect 181363 110866 181683 110898
rect 181794 111454 182414 146898
rect 185514 151174 186134 177223
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 184836 115174 185156 115206
rect 184836 114938 184878 115174
rect 185114 114938 185156 115174
rect 184836 114854 185156 114938
rect 184836 114618 184878 114854
rect 185114 114618 185156 114854
rect 184836 114586 185156 114618
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 189234 154894 189854 170068
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 115001 189854 118338
rect 192954 158614 193574 177223
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 191782 115174 192102 115206
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 171834 101258 171866 101494
rect 172102 101258 172186 101494
rect 172422 101258 172454 101494
rect 171834 101174 172454 101258
rect 171834 100938 171866 101174
rect 172102 100938 172186 101174
rect 172422 100938 172454 101174
rect 170075 98972 170141 98973
rect 170075 98908 170076 98972
rect 170140 98908 170141 98972
rect 170075 98907 170141 98908
rect 170078 57221 170138 98907
rect 170259 73812 170325 73813
rect 170259 73748 170260 73812
rect 170324 73748 170325 73812
rect 170259 73747 170325 73748
rect 170262 69733 170322 73747
rect 170259 69732 170325 69733
rect 170259 69668 170260 69732
rect 170324 69668 170325 69732
rect 170259 69667 170325 69668
rect 171834 65494 172454 100938
rect 177890 79174 178210 79206
rect 177890 78938 177932 79174
rect 178168 78938 178210 79174
rect 177890 78854 178210 78938
rect 177890 78618 177932 78854
rect 178168 78618 178210 78854
rect 177890 78586 178210 78618
rect 174417 75454 174737 75486
rect 174417 75218 174459 75454
rect 174695 75218 174737 75454
rect 174417 75134 174737 75218
rect 174417 74898 174459 75134
rect 174695 74898 174737 75134
rect 174417 74866 174737 74898
rect 181363 75454 181683 75486
rect 181363 75218 181405 75454
rect 181641 75218 181683 75454
rect 181363 75134 181683 75218
rect 181363 74898 181405 75134
rect 181641 74898 181683 75134
rect 181363 74866 181683 74898
rect 181794 75454 182414 110898
rect 184836 79174 185156 79206
rect 184836 78938 184878 79174
rect 185114 78938 185156 79174
rect 184836 78854 185156 78938
rect 184836 78618 184878 78854
rect 185114 78618 185156 78854
rect 184836 78586 185156 78618
rect 185514 79174 186134 114618
rect 191782 114938 191824 115174
rect 192060 114938 192102 115174
rect 191782 114854 192102 114938
rect 191782 114618 191824 114854
rect 192060 114618 192102 114854
rect 191782 114586 192102 114618
rect 188309 111454 188629 111486
rect 188309 111218 188351 111454
rect 188587 111218 188629 111454
rect 188309 111134 188629 111218
rect 188309 110898 188351 111134
rect 188587 110898 188629 111134
rect 188309 110866 188629 110898
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 171834 65258 171866 65494
rect 172102 65258 172186 65494
rect 172422 65258 172454 65494
rect 171834 65174 172454 65258
rect 171834 64938 171866 65174
rect 172102 64938 172186 65174
rect 172422 64938 172454 65174
rect 170075 57220 170141 57221
rect 170075 57156 170076 57220
rect 170140 57156 170141 57220
rect 170075 57155 170141 57156
rect 169891 40628 169957 40629
rect 169891 40564 169892 40628
rect 169956 40564 169957 40628
rect 169891 40563 169957 40564
rect 171834 29494 172454 64938
rect 171834 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 172454 29494
rect 171834 29174 172454 29258
rect 171834 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 172454 29174
rect 169523 19956 169589 19957
rect 169523 19892 169524 19956
rect 169588 19892 169589 19956
rect 169523 19891 169589 19892
rect 168114 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 168734 -6106
rect 168114 -6426 168734 -6342
rect 168114 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 168734 -6426
rect 168114 -7654 168734 -6662
rect 171834 -7066 172454 28938
rect 171834 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 172454 -7066
rect 171834 -7386 172454 -7302
rect 171834 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 172454 -7386
rect 171834 -7654 172454 -7622
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 185514 43174 186134 78618
rect 189234 82894 189854 92591
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 188309 75454 188629 75486
rect 188309 75218 188351 75454
rect 188587 75218 188629 75454
rect 188309 75134 188629 75218
rect 188309 74898 188351 75134
rect 188587 74898 188629 75134
rect 188309 74866 188629 74898
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -1306 186134 6618
rect 185514 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 186134 -1306
rect 185514 -1626 186134 -1542
rect 185514 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 186134 -1626
rect 185514 -7654 186134 -1862
rect 189234 46894 189854 82338
rect 192954 86614 193574 122058
rect 196674 162334 197294 177223
rect 199331 168332 199397 168333
rect 199331 168268 199332 168332
rect 199396 168268 199397 168332
rect 199331 168267 199397 168268
rect 196674 162098 196706 162334
rect 196942 162098 197026 162334
rect 197262 162098 197294 162334
rect 196674 162014 197294 162098
rect 196674 161778 196706 162014
rect 196942 161778 197026 162014
rect 197262 161778 197294 162014
rect 196674 126334 197294 161778
rect 196674 126098 196706 126334
rect 196942 126098 197026 126334
rect 197262 126098 197294 126334
rect 196674 126014 197294 126098
rect 196674 125778 196706 126014
rect 196942 125778 197026 126014
rect 197262 125778 197294 126014
rect 195255 111454 195575 111486
rect 195255 111218 195297 111454
rect 195533 111218 195575 111454
rect 195255 111134 195575 111218
rect 195255 110898 195297 111134
rect 195533 110898 195575 111134
rect 195255 110866 195575 110898
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 191782 79174 192102 79206
rect 191782 78938 191824 79174
rect 192060 78938 192102 79174
rect 191782 78854 192102 78938
rect 191782 78618 191824 78854
rect 192060 78618 192102 78854
rect 191782 78586 192102 78618
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -2266 189854 10338
rect 189234 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 189854 -2266
rect 189234 -2586 189854 -2502
rect 189234 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 189854 -2586
rect 189234 -7654 189854 -2822
rect 192954 50614 193574 86058
rect 196674 90334 197294 125778
rect 198728 115174 199048 115206
rect 198728 114938 198770 115174
rect 199006 114938 199048 115174
rect 198728 114854 199048 114938
rect 198728 114618 198770 114854
rect 199006 114618 199048 114854
rect 198728 114586 199048 114618
rect 199334 113250 199394 168267
rect 200394 166054 201014 177223
rect 200394 165818 200426 166054
rect 200662 165818 200746 166054
rect 200982 165818 201014 166054
rect 200394 165734 201014 165818
rect 200394 165498 200426 165734
rect 200662 165498 200746 165734
rect 200982 165498 201014 165734
rect 200394 130054 201014 165498
rect 200394 129818 200426 130054
rect 200662 129818 200746 130054
rect 200982 129818 201014 130054
rect 200394 129734 201014 129818
rect 200394 129498 200426 129734
rect 200662 129498 200746 129734
rect 200982 129498 201014 129734
rect 199515 124268 199581 124269
rect 199515 124204 199516 124268
rect 199580 124204 199581 124268
rect 199515 124203 199581 124204
rect 199518 116381 199578 124203
rect 200067 119372 200133 119373
rect 200067 119370 200068 119372
rect 199702 119310 200068 119370
rect 199702 119101 199762 119310
rect 200067 119308 200068 119310
rect 200132 119308 200133 119372
rect 200067 119307 200133 119308
rect 199699 119100 199765 119101
rect 199699 119036 199700 119100
rect 199764 119036 199765 119100
rect 199699 119035 199765 119036
rect 200067 118692 200133 118693
rect 200067 118690 200068 118692
rect 199702 118630 200068 118690
rect 199702 118421 199762 118630
rect 200067 118628 200068 118630
rect 200132 118628 200133 118692
rect 200067 118627 200133 118628
rect 199699 118420 199765 118421
rect 199699 118356 199700 118420
rect 199764 118356 199765 118420
rect 199699 118355 199765 118356
rect 200067 118012 200133 118013
rect 200067 118010 200068 118012
rect 199702 117950 200068 118010
rect 199702 117741 199762 117950
rect 200067 117948 200068 117950
rect 200132 117948 200133 118012
rect 200067 117947 200133 117948
rect 199699 117740 199765 117741
rect 199699 117676 199700 117740
rect 199764 117676 199765 117740
rect 199699 117675 199765 117676
rect 200067 117332 200133 117333
rect 200067 117330 200068 117332
rect 199702 117270 200068 117330
rect 199702 117061 199762 117270
rect 200067 117268 200068 117270
rect 200132 117268 200133 117332
rect 200067 117267 200133 117268
rect 199699 117060 199765 117061
rect 199699 116996 199700 117060
rect 199764 116996 199765 117060
rect 199699 116995 199765 116996
rect 199515 116380 199581 116381
rect 199515 116316 199516 116380
rect 199580 116316 199581 116380
rect 199515 116315 199581 116316
rect 200067 115972 200133 115973
rect 200067 115970 200068 115972
rect 199702 115910 200068 115970
rect 199702 115701 199762 115910
rect 200067 115908 200068 115910
rect 200132 115908 200133 115972
rect 200067 115907 200133 115908
rect 199699 115700 199765 115701
rect 199699 115636 199700 115700
rect 199764 115636 199765 115700
rect 199699 115635 199765 115636
rect 200067 115292 200133 115293
rect 200067 115290 200068 115292
rect 199702 115230 200068 115290
rect 199702 115021 199762 115230
rect 200067 115228 200068 115230
rect 200132 115228 200133 115292
rect 200067 115227 200133 115228
rect 199699 115020 199765 115021
rect 199699 114956 199700 115020
rect 199764 114956 199765 115020
rect 199699 114955 199765 114956
rect 200067 114612 200133 114613
rect 200067 114610 200068 114612
rect 199702 114550 200068 114610
rect 199702 113661 199762 114550
rect 200067 114548 200068 114550
rect 200132 114548 200133 114612
rect 200067 114547 200133 114548
rect 199699 113660 199765 113661
rect 199699 113596 199700 113660
rect 199764 113596 199765 113660
rect 199699 113595 199765 113596
rect 200067 113252 200133 113253
rect 200067 113250 200068 113252
rect 199334 113190 200068 113250
rect 200067 113188 200068 113190
rect 200132 113188 200133 113252
rect 200067 113187 200133 113188
rect 199699 112844 199765 112845
rect 199699 112780 199700 112844
rect 199764 112780 199765 112844
rect 199699 112779 199765 112780
rect 199702 112570 199762 112779
rect 200067 112572 200133 112573
rect 200067 112570 200068 112572
rect 199702 112510 200068 112570
rect 200067 112508 200068 112510
rect 200132 112508 200133 112572
rect 200067 112507 200133 112508
rect 199699 112164 199765 112165
rect 199699 112100 199700 112164
rect 199764 112100 199765 112164
rect 199699 112099 199765 112100
rect 199702 111890 199762 112099
rect 200067 111892 200133 111893
rect 200067 111890 200068 111892
rect 199702 111830 200068 111890
rect 200067 111828 200068 111830
rect 200132 111828 200133 111892
rect 200067 111827 200133 111828
rect 199699 111484 199765 111485
rect 199699 111420 199700 111484
rect 199764 111420 199765 111484
rect 199699 111419 199765 111420
rect 199702 111210 199762 111419
rect 200067 111212 200133 111213
rect 200067 111210 200068 111212
rect 199702 111150 200068 111210
rect 200067 111148 200068 111150
rect 200132 111148 200133 111212
rect 200067 111147 200133 111148
rect 199699 110804 199765 110805
rect 199699 110740 199700 110804
rect 199764 110740 199765 110804
rect 199699 110739 199765 110740
rect 199702 110530 199762 110739
rect 200067 110532 200133 110533
rect 200067 110530 200068 110532
rect 199702 110470 200068 110530
rect 200067 110468 200068 110470
rect 200132 110468 200133 110532
rect 200067 110467 200133 110468
rect 199699 110124 199765 110125
rect 199699 110060 199700 110124
rect 199764 110060 199765 110124
rect 199699 110059 199765 110060
rect 199702 109850 199762 110059
rect 200067 109852 200133 109853
rect 200067 109850 200068 109852
rect 199702 109790 200068 109850
rect 200067 109788 200068 109790
rect 200132 109788 200133 109852
rect 200067 109787 200133 109788
rect 199699 109444 199765 109445
rect 199699 109380 199700 109444
rect 199764 109380 199765 109444
rect 199699 109379 199765 109380
rect 199702 109170 199762 109379
rect 200067 109172 200133 109173
rect 200067 109170 200068 109172
rect 199702 109110 200068 109170
rect 200067 109108 200068 109110
rect 200132 109108 200133 109172
rect 200067 109107 200133 109108
rect 200067 108492 200133 108493
rect 200067 108490 200068 108492
rect 199702 108430 200068 108490
rect 199702 108221 199762 108430
rect 200067 108428 200068 108430
rect 200132 108428 200133 108492
rect 200067 108427 200133 108428
rect 199699 108220 199765 108221
rect 199699 108156 199700 108220
rect 199764 108156 199765 108220
rect 199699 108155 199765 108156
rect 199699 107404 199765 107405
rect 199699 107340 199700 107404
rect 199764 107340 199765 107404
rect 199699 107339 199765 107340
rect 199702 107130 199762 107339
rect 200067 107132 200133 107133
rect 200067 107130 200068 107132
rect 199702 107070 200068 107130
rect 200067 107068 200068 107070
rect 200132 107068 200133 107132
rect 200067 107067 200133 107068
rect 199699 106724 199765 106725
rect 199699 106660 199700 106724
rect 199764 106660 199765 106724
rect 199699 106659 199765 106660
rect 199702 106450 199762 106659
rect 200067 106452 200133 106453
rect 200067 106450 200068 106452
rect 199702 106390 200068 106450
rect 200067 106388 200068 106390
rect 200132 106388 200133 106452
rect 200067 106387 200133 106388
rect 199515 106044 199581 106045
rect 199515 105980 199516 106044
rect 199580 105980 199581 106044
rect 199515 105979 199581 105980
rect 199518 105090 199578 105979
rect 200067 105772 200133 105773
rect 200067 105770 200068 105772
rect 199702 105710 200068 105770
rect 199702 105501 199762 105710
rect 200067 105708 200068 105710
rect 200132 105708 200133 105772
rect 200067 105707 200133 105708
rect 199699 105500 199765 105501
rect 199699 105436 199700 105500
rect 199764 105436 199765 105500
rect 199699 105435 199765 105436
rect 200067 105092 200133 105093
rect 200067 105090 200068 105092
rect 199518 105030 200068 105090
rect 200067 105028 200068 105030
rect 200132 105028 200133 105092
rect 200067 105027 200133 105028
rect 199515 104684 199581 104685
rect 199515 104620 199516 104684
rect 199580 104620 199581 104684
rect 199515 104619 199581 104620
rect 199518 103730 199578 104619
rect 200067 104412 200133 104413
rect 200067 104410 200068 104412
rect 199702 104350 200068 104410
rect 199702 104141 199762 104350
rect 200067 104348 200068 104350
rect 200132 104348 200133 104412
rect 200067 104347 200133 104348
rect 199699 104140 199765 104141
rect 199699 104076 199700 104140
rect 199764 104076 199765 104140
rect 199699 104075 199765 104076
rect 200067 103732 200133 103733
rect 200067 103730 200068 103732
rect 199518 103670 200068 103730
rect 200067 103668 200068 103670
rect 200132 103668 200133 103732
rect 200067 103667 200133 103668
rect 200067 103052 200133 103053
rect 200067 103050 200068 103052
rect 199702 102990 200068 103050
rect 199702 102781 199762 102990
rect 200067 102988 200068 102990
rect 200132 102988 200133 103052
rect 200067 102987 200133 102988
rect 199699 102780 199765 102781
rect 199699 102716 199700 102780
rect 199764 102716 199765 102780
rect 199699 102715 199765 102716
rect 199699 101964 199765 101965
rect 199699 101900 199700 101964
rect 199764 101900 199765 101964
rect 199699 101899 199765 101900
rect 199702 101690 199762 101899
rect 200067 101692 200133 101693
rect 200067 101690 200068 101692
rect 199702 101630 200068 101690
rect 200067 101628 200068 101630
rect 200132 101628 200133 101692
rect 200067 101627 200133 101628
rect 199699 101284 199765 101285
rect 199699 101220 199700 101284
rect 199764 101220 199765 101284
rect 199699 101219 199765 101220
rect 199702 101010 199762 101219
rect 200067 101012 200133 101013
rect 200067 101010 200068 101012
rect 199702 100950 200068 101010
rect 200067 100948 200068 100950
rect 200132 100948 200133 101012
rect 200067 100947 200133 100948
rect 199699 100604 199765 100605
rect 199699 100540 199700 100604
rect 199764 100540 199765 100604
rect 199699 100539 199765 100540
rect 199702 100330 199762 100539
rect 200067 100332 200133 100333
rect 200067 100330 200068 100332
rect 199702 100270 200068 100330
rect 200067 100268 200068 100270
rect 200132 100268 200133 100332
rect 200067 100267 200133 100268
rect 199699 99924 199765 99925
rect 199699 99860 199700 99924
rect 199764 99860 199765 99924
rect 199699 99859 199765 99860
rect 199702 99650 199762 99859
rect 200067 99652 200133 99653
rect 200067 99650 200068 99652
rect 199702 99590 200068 99650
rect 200067 99588 200068 99590
rect 200132 99588 200133 99652
rect 200067 99587 200133 99588
rect 199699 99244 199765 99245
rect 199699 99180 199700 99244
rect 199764 99180 199765 99244
rect 199699 99179 199765 99180
rect 199702 98970 199762 99179
rect 200067 98972 200133 98973
rect 200067 98970 200068 98972
rect 199702 98910 200068 98970
rect 200067 98908 200068 98910
rect 200132 98908 200133 98972
rect 200067 98907 200133 98908
rect 199699 98564 199765 98565
rect 199699 98500 199700 98564
rect 199764 98500 199765 98564
rect 199699 98499 199765 98500
rect 199702 98290 199762 98499
rect 200067 98292 200133 98293
rect 200067 98290 200068 98292
rect 199702 98230 200068 98290
rect 200067 98228 200068 98230
rect 200132 98228 200133 98292
rect 200067 98227 200133 98228
rect 200067 97612 200133 97613
rect 200067 97610 200068 97612
rect 199702 97550 200068 97610
rect 199702 97341 199762 97550
rect 200067 97548 200068 97550
rect 200132 97548 200133 97612
rect 200067 97547 200133 97548
rect 199699 97340 199765 97341
rect 199699 97276 199700 97340
rect 199764 97276 199765 97340
rect 199699 97275 199765 97276
rect 200067 96932 200133 96933
rect 200067 96930 200068 96932
rect 199702 96870 200068 96930
rect 199702 96661 199762 96870
rect 200067 96868 200068 96870
rect 200132 96868 200133 96932
rect 200067 96867 200133 96868
rect 199699 96660 199765 96661
rect 199699 96596 199700 96660
rect 199764 96596 199765 96660
rect 199699 96595 199765 96596
rect 200067 96252 200133 96253
rect 200067 96250 200068 96252
rect 199702 96190 200068 96250
rect 199702 95981 199762 96190
rect 200067 96188 200068 96190
rect 200132 96188 200133 96252
rect 200067 96187 200133 96188
rect 199699 95980 199765 95981
rect 199699 95916 199700 95980
rect 199764 95916 199765 95980
rect 199699 95915 199765 95916
rect 200067 95572 200133 95573
rect 200067 95570 200068 95572
rect 199702 95510 200068 95570
rect 199702 95301 199762 95510
rect 200067 95508 200068 95510
rect 200132 95508 200133 95572
rect 200067 95507 200133 95508
rect 199699 95300 199765 95301
rect 199699 95236 199700 95300
rect 199764 95236 199765 95300
rect 199699 95235 199765 95236
rect 200067 94892 200133 94893
rect 200067 94890 200068 94892
rect 199702 94830 200068 94890
rect 199702 94621 199762 94830
rect 200067 94828 200068 94830
rect 200132 94828 200133 94892
rect 200067 94827 200133 94828
rect 199699 94620 199765 94621
rect 199699 94556 199700 94620
rect 199764 94556 199765 94620
rect 199699 94555 199765 94556
rect 200067 94212 200133 94213
rect 200067 94210 200068 94212
rect 199702 94150 200068 94210
rect 199702 93941 199762 94150
rect 200067 94148 200068 94150
rect 200132 94148 200133 94212
rect 200067 94147 200133 94148
rect 200394 94054 201014 129498
rect 204114 169774 204734 177223
rect 204114 169538 204146 169774
rect 204382 169538 204466 169774
rect 204702 169538 204734 169774
rect 204114 169454 204734 169538
rect 204114 169218 204146 169454
rect 204382 169218 204466 169454
rect 204702 169218 204734 169454
rect 204114 133774 204734 169218
rect 204114 133538 204146 133774
rect 204382 133538 204466 133774
rect 204702 133538 204734 133774
rect 204114 133454 204734 133538
rect 204114 133218 204146 133454
rect 204382 133218 204466 133454
rect 204702 133218 204734 133454
rect 201539 101012 201605 101013
rect 201539 100948 201540 101012
rect 201604 100948 201605 101012
rect 201539 100947 201605 100948
rect 199699 93940 199765 93941
rect 199699 93876 199700 93940
rect 199764 93876 199765 93940
rect 199699 93875 199765 93876
rect 200394 93818 200426 94054
rect 200662 93818 200746 94054
rect 200982 93818 201014 94054
rect 200394 93734 201014 93818
rect 200394 93498 200426 93734
rect 200662 93498 200746 93734
rect 200982 93498 201014 93734
rect 199699 93124 199765 93125
rect 199699 93060 199700 93124
rect 199764 93060 199765 93124
rect 199699 93059 199765 93060
rect 199702 92850 199762 93059
rect 200067 92852 200133 92853
rect 200067 92850 200068 92852
rect 199702 92790 200068 92850
rect 200067 92788 200068 92790
rect 200132 92788 200133 92852
rect 200067 92787 200133 92788
rect 200067 92172 200133 92173
rect 200067 92170 200068 92172
rect 199702 92110 200068 92170
rect 199702 91901 199762 92110
rect 200067 92108 200068 92110
rect 200132 92108 200133 92172
rect 200067 92107 200133 92108
rect 199699 91900 199765 91901
rect 199699 91836 199700 91900
rect 199764 91836 199765 91900
rect 199699 91835 199765 91836
rect 200067 91492 200133 91493
rect 200067 91490 200068 91492
rect 199702 91430 200068 91490
rect 199702 91221 199762 91430
rect 200067 91428 200068 91430
rect 200132 91428 200133 91492
rect 200067 91427 200133 91428
rect 199699 91220 199765 91221
rect 199699 91156 199700 91220
rect 199764 91156 199765 91220
rect 199699 91155 199765 91156
rect 200067 90812 200133 90813
rect 200067 90810 200068 90812
rect 199702 90750 200068 90810
rect 199702 90541 199762 90750
rect 200067 90748 200068 90750
rect 200132 90748 200133 90812
rect 200067 90747 200133 90748
rect 199699 90540 199765 90541
rect 199699 90476 199700 90540
rect 199764 90476 199765 90540
rect 199699 90475 199765 90476
rect 196674 90098 196706 90334
rect 196942 90098 197026 90334
rect 197262 90098 197294 90334
rect 200067 90132 200133 90133
rect 200067 90130 200068 90132
rect 196674 90014 197294 90098
rect 196674 89778 196706 90014
rect 196942 89778 197026 90014
rect 197262 89778 197294 90014
rect 199702 90070 200068 90130
rect 199702 89861 199762 90070
rect 200067 90068 200068 90070
rect 200132 90068 200133 90132
rect 200067 90067 200133 90068
rect 199699 89860 199765 89861
rect 199699 89796 199700 89860
rect 199764 89796 199765 89860
rect 199699 89795 199765 89796
rect 195255 75454 195575 75486
rect 195255 75218 195297 75454
rect 195533 75218 195575 75454
rect 195255 75134 195575 75218
rect 195255 74898 195297 75134
rect 195533 74898 195575 75134
rect 195255 74866 195575 74898
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 192954 -3226 193574 14058
rect 192954 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 193574 -3226
rect 192954 -3546 193574 -3462
rect 192954 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 193574 -3546
rect 192954 -7654 193574 -3782
rect 196674 54334 197294 89778
rect 200067 89452 200133 89453
rect 200067 89450 200068 89452
rect 199702 89390 200068 89450
rect 199702 89181 199762 89390
rect 200067 89388 200068 89390
rect 200132 89388 200133 89452
rect 200067 89387 200133 89388
rect 199699 89180 199765 89181
rect 199699 89116 199700 89180
rect 199764 89116 199765 89180
rect 199699 89115 199765 89116
rect 200067 88772 200133 88773
rect 200067 88770 200068 88772
rect 199702 88710 200068 88770
rect 199702 88501 199762 88710
rect 200067 88708 200068 88710
rect 200132 88708 200133 88772
rect 200067 88707 200133 88708
rect 199699 88500 199765 88501
rect 199699 88436 199700 88500
rect 199764 88436 199765 88500
rect 199699 88435 199765 88436
rect 200067 88092 200133 88093
rect 200067 88090 200068 88092
rect 199702 88030 200068 88090
rect 199702 87821 199762 88030
rect 200067 88028 200068 88030
rect 200132 88028 200133 88092
rect 200067 88027 200133 88028
rect 199699 87820 199765 87821
rect 199699 87756 199700 87820
rect 199764 87756 199765 87820
rect 199699 87755 199765 87756
rect 200067 86732 200133 86733
rect 200067 86730 200068 86732
rect 199702 86670 200068 86730
rect 199702 86461 199762 86670
rect 200067 86668 200068 86670
rect 200132 86668 200133 86732
rect 200067 86667 200133 86668
rect 199699 86460 199765 86461
rect 199699 86396 199700 86460
rect 199764 86396 199765 86460
rect 199699 86395 199765 86396
rect 200067 86052 200133 86053
rect 200067 86050 200068 86052
rect 199150 85990 200068 86050
rect 199150 80070 199210 85990
rect 200067 85988 200068 85990
rect 200132 85988 200133 86052
rect 200067 85987 200133 85988
rect 199699 85644 199765 85645
rect 199699 85580 199700 85644
rect 199764 85580 199765 85644
rect 199699 85579 199765 85580
rect 200067 85644 200133 85645
rect 200067 85580 200068 85644
rect 200132 85580 200133 85644
rect 200067 85579 200133 85580
rect 199702 85370 199762 85579
rect 200070 85370 200130 85579
rect 199702 85310 200130 85370
rect 199699 84964 199765 84965
rect 199699 84900 199700 84964
rect 199764 84900 199765 84964
rect 199699 84899 199765 84900
rect 199702 84690 199762 84899
rect 200067 84828 200133 84829
rect 200067 84764 200068 84828
rect 200132 84764 200133 84828
rect 200067 84763 200133 84764
rect 200070 84690 200130 84763
rect 199702 84630 200130 84690
rect 199699 84284 199765 84285
rect 199699 84220 199700 84284
rect 199764 84220 199765 84284
rect 199699 84219 199765 84220
rect 200067 84284 200133 84285
rect 200067 84220 200068 84284
rect 200132 84220 200133 84284
rect 200067 84219 200133 84220
rect 199702 84010 199762 84219
rect 200070 84010 200130 84219
rect 199702 83950 200130 84010
rect 199331 83604 199397 83605
rect 199331 83540 199332 83604
rect 199396 83540 199397 83604
rect 199331 83539 199397 83540
rect 199334 82650 199394 83539
rect 200067 83332 200133 83333
rect 200067 83330 200068 83332
rect 199702 83270 200068 83330
rect 199702 83061 199762 83270
rect 200067 83268 200068 83270
rect 200132 83268 200133 83332
rect 200067 83267 200133 83268
rect 199699 83060 199765 83061
rect 199699 82996 199700 83060
rect 199764 82996 199765 83060
rect 199699 82995 199765 82996
rect 200067 82924 200133 82925
rect 200067 82860 200068 82924
rect 200132 82860 200133 82924
rect 200067 82859 200133 82860
rect 200070 82650 200130 82859
rect 199334 82590 200130 82650
rect 199699 82244 199765 82245
rect 199699 82180 199700 82244
rect 199764 82180 199765 82244
rect 199699 82179 199765 82180
rect 199702 81970 199762 82179
rect 200067 81972 200133 81973
rect 200067 81970 200068 81972
rect 199702 81910 200068 81970
rect 200067 81908 200068 81910
rect 200132 81908 200133 81972
rect 200067 81907 200133 81908
rect 199699 80884 199765 80885
rect 199699 80820 199700 80884
rect 199764 80820 199765 80884
rect 199699 80819 199765 80820
rect 199702 80610 199762 80819
rect 200067 80612 200133 80613
rect 200067 80610 200068 80612
rect 199702 80550 200068 80610
rect 200067 80548 200068 80550
rect 200132 80548 200133 80612
rect 200067 80547 200133 80548
rect 199699 80204 199765 80205
rect 199699 80140 199700 80204
rect 199764 80140 199765 80204
rect 199699 80139 199765 80140
rect 199702 80070 199762 80139
rect 199150 80010 199578 80070
rect 199702 80069 200130 80070
rect 199702 80068 200133 80069
rect 199702 80010 200068 80068
rect 198728 79174 199048 79206
rect 198728 78938 198770 79174
rect 199006 78938 199048 79174
rect 198728 78854 199048 78938
rect 198728 78618 198770 78854
rect 199006 78618 199048 78854
rect 198728 78586 199048 78618
rect 199331 78164 199397 78165
rect 199331 78100 199332 78164
rect 199396 78100 199397 78164
rect 199331 78099 199397 78100
rect 199334 75170 199394 78099
rect 199518 75850 199578 80010
rect 200067 80004 200068 80010
rect 200132 80004 200133 80068
rect 200067 80003 200133 80004
rect 199699 79524 199765 79525
rect 199699 79460 199700 79524
rect 199764 79460 199765 79524
rect 199699 79459 199765 79460
rect 199702 79250 199762 79459
rect 200067 79252 200133 79253
rect 200067 79250 200068 79252
rect 199702 79190 200068 79250
rect 200067 79188 200068 79190
rect 200132 79188 200133 79252
rect 200067 79187 200133 79188
rect 199699 78844 199765 78845
rect 199699 78780 199700 78844
rect 199764 78780 199765 78844
rect 199699 78779 199765 78780
rect 199702 78570 199762 78779
rect 200067 78708 200133 78709
rect 200067 78644 200068 78708
rect 200132 78644 200133 78708
rect 200067 78643 200133 78644
rect 200070 78570 200130 78643
rect 199702 78510 200130 78570
rect 199699 77484 199765 77485
rect 199699 77420 199700 77484
rect 199764 77420 199765 77484
rect 199699 77419 199765 77420
rect 199702 77210 199762 77419
rect 200067 77348 200133 77349
rect 200067 77284 200068 77348
rect 200132 77284 200133 77348
rect 200067 77283 200133 77284
rect 200070 77210 200130 77283
rect 199702 77150 200130 77210
rect 199699 76804 199765 76805
rect 199699 76740 199700 76804
rect 199764 76740 199765 76804
rect 199699 76739 199765 76740
rect 199702 76530 199762 76739
rect 200067 76532 200133 76533
rect 200067 76530 200068 76532
rect 199702 76470 200068 76530
rect 200067 76468 200068 76470
rect 200132 76468 200133 76532
rect 200067 76467 200133 76468
rect 199518 75790 200314 75850
rect 199699 75444 199765 75445
rect 199699 75380 199700 75444
rect 199764 75380 199765 75444
rect 199699 75379 199765 75380
rect 199150 75110 199394 75170
rect 199702 75170 199762 75379
rect 200067 75172 200133 75173
rect 200067 75170 200068 75172
rect 199702 75110 200068 75170
rect 199150 69325 199210 75110
rect 200067 75108 200068 75110
rect 200132 75108 200133 75172
rect 200067 75107 200133 75108
rect 199331 74764 199397 74765
rect 199331 74700 199332 74764
rect 199396 74762 199397 74764
rect 200067 74764 200133 74765
rect 200067 74762 200068 74764
rect 199396 74702 200068 74762
rect 199396 74700 199397 74702
rect 199331 74699 199397 74700
rect 200067 74700 200068 74702
rect 200132 74700 200133 74764
rect 200067 74699 200133 74700
rect 199334 69461 199394 74699
rect 199699 74084 199765 74085
rect 199699 74020 199700 74084
rect 199764 74020 199765 74084
rect 199699 74019 199765 74020
rect 199702 73810 199762 74019
rect 200067 73812 200133 73813
rect 200067 73810 200068 73812
rect 199702 73750 200068 73810
rect 200067 73748 200068 73750
rect 200132 73748 200133 73812
rect 200067 73747 200133 73748
rect 199699 73404 199765 73405
rect 199699 73340 199700 73404
rect 199764 73340 199765 73404
rect 199699 73339 199765 73340
rect 199702 73130 199762 73339
rect 200067 73268 200133 73269
rect 200067 73204 200068 73268
rect 200132 73204 200133 73268
rect 200067 73203 200133 73204
rect 200070 73130 200130 73203
rect 199702 73070 200130 73130
rect 199699 72724 199765 72725
rect 199699 72660 199700 72724
rect 199764 72660 199765 72724
rect 199699 72659 199765 72660
rect 199702 72450 199762 72659
rect 200067 72452 200133 72453
rect 200067 72450 200068 72452
rect 199702 72390 200068 72450
rect 200067 72388 200068 72390
rect 200132 72388 200133 72452
rect 200067 72387 200133 72388
rect 199699 72044 199765 72045
rect 199699 71980 199700 72044
rect 199764 71980 199765 72044
rect 199699 71979 199765 71980
rect 199702 71770 199762 71979
rect 200067 71908 200133 71909
rect 200067 71844 200068 71908
rect 200132 71844 200133 71908
rect 200067 71843 200133 71844
rect 200070 71770 200130 71843
rect 199702 71710 200130 71770
rect 199331 69460 199397 69461
rect 199331 69396 199332 69460
rect 199396 69396 199397 69460
rect 199331 69395 199397 69396
rect 199147 69324 199213 69325
rect 199147 69260 199148 69324
rect 199212 69260 199213 69324
rect 199147 69259 199213 69260
rect 200067 68916 200133 68917
rect 200067 68852 200068 68916
rect 200132 68914 200133 68916
rect 200254 68914 200314 75790
rect 200132 68854 200314 68914
rect 200132 68852 200133 68854
rect 200067 68851 200133 68852
rect 196674 54098 196706 54334
rect 196942 54098 197026 54334
rect 197262 54098 197294 54334
rect 196674 54014 197294 54098
rect 196674 53778 196706 54014
rect 196942 53778 197026 54014
rect 197262 53778 197294 54014
rect 196674 18334 197294 53778
rect 196674 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 197294 18334
rect 196674 18014 197294 18098
rect 196674 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 197294 18014
rect 196674 -4186 197294 17778
rect 196674 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 197294 -4186
rect 196674 -4506 197294 -4422
rect 196674 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 197294 -4506
rect 196674 -7654 197294 -4742
rect 200394 58054 201014 93498
rect 201542 67285 201602 100947
rect 204114 97774 204734 133218
rect 204114 97538 204146 97774
rect 204382 97538 204466 97774
rect 204702 97538 204734 97774
rect 204114 97454 204734 97538
rect 204114 97218 204146 97454
rect 204382 97218 204466 97454
rect 204702 97218 204734 97454
rect 201723 91492 201789 91493
rect 201723 91428 201724 91492
rect 201788 91428 201789 91492
rect 201723 91427 201789 91428
rect 201726 69597 201786 91427
rect 201723 69596 201789 69597
rect 201723 69532 201724 69596
rect 201788 69532 201789 69596
rect 201723 69531 201789 69532
rect 201539 67284 201605 67285
rect 201539 67220 201540 67284
rect 201604 67220 201605 67284
rect 201539 67219 201605 67220
rect 200394 57818 200426 58054
rect 200662 57818 200746 58054
rect 200982 57818 201014 58054
rect 200394 57734 201014 57818
rect 200394 57498 200426 57734
rect 200662 57498 200746 57734
rect 200982 57498 201014 57734
rect 200394 22054 201014 57498
rect 200394 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 201014 22054
rect 200394 21734 201014 21818
rect 200394 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 201014 21734
rect 200394 -5146 201014 21498
rect 200394 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 201014 -5146
rect 200394 -5466 201014 -5382
rect 200394 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 201014 -5466
rect 200394 -7654 201014 -5702
rect 204114 61774 204734 97218
rect 204114 61538 204146 61774
rect 204382 61538 204466 61774
rect 204702 61538 204734 61774
rect 204114 61454 204734 61538
rect 204114 61218 204146 61454
rect 204382 61218 204466 61454
rect 204702 61218 204734 61454
rect 204114 25774 204734 61218
rect 204114 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 204734 25774
rect 204114 25454 204734 25538
rect 204114 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 204734 25454
rect 204114 -6106 204734 25218
rect 204114 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 204734 -6106
rect 204114 -6426 204734 -6342
rect 204114 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 204734 -6426
rect 204114 -7654 204734 -6662
rect 207834 173494 208454 177223
rect 207834 173258 207866 173494
rect 208102 173258 208186 173494
rect 208422 173258 208454 173494
rect 207834 173174 208454 173258
rect 207834 172938 207866 173174
rect 208102 172938 208186 173174
rect 208422 172938 208454 173174
rect 207834 137494 208454 172938
rect 207834 137258 207866 137494
rect 208102 137258 208186 137494
rect 208422 137258 208454 137494
rect 207834 137174 208454 137258
rect 207834 136938 207866 137174
rect 208102 136938 208186 137174
rect 208422 136938 208454 137174
rect 207834 101494 208454 136938
rect 207834 101258 207866 101494
rect 208102 101258 208186 101494
rect 208422 101258 208454 101494
rect 207834 101174 208454 101258
rect 207834 100938 207866 101174
rect 208102 100938 208186 101174
rect 208422 100938 208454 101174
rect 207834 65494 208454 100938
rect 207834 65258 207866 65494
rect 208102 65258 208186 65494
rect 208422 65258 208454 65494
rect 207834 65174 208454 65258
rect 207834 64938 207866 65174
rect 208102 64938 208186 65174
rect 208422 64938 208454 65174
rect 207834 29494 208454 64938
rect 207834 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 208454 29494
rect 207834 29174 208454 29258
rect 207834 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 208454 29174
rect 207834 -7066 208454 28938
rect 207834 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 208454 -7066
rect 207834 -7386 208454 -7302
rect 207834 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 208454 -7386
rect 207834 -7654 208454 -7622
rect 217794 147454 218414 177223
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 221514 151174 222134 186618
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 115174 222134 150618
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -1306 222134 6618
rect 221514 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 222134 -1306
rect 221514 -1626 222134 -1542
rect 221514 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 222134 -1626
rect 221514 -7654 222134 -1862
rect 225234 706758 225854 711590
rect 225234 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 225854 706758
rect 225234 706438 225854 706522
rect 225234 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 225854 706438
rect 225234 694894 225854 706202
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 262894 225854 298338
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 226894 225854 262338
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 154894 225854 190338
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 118894 225854 154338
rect 225234 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 225854 118894
rect 225234 118574 225854 118658
rect 225234 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 225854 118574
rect 225234 82894 225854 118338
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -2266 225854 10338
rect 225234 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 225854 -2266
rect 225234 -2586 225854 -2502
rect 225234 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 225854 -2586
rect 225234 -7654 225854 -2822
rect 228954 707718 229574 711590
rect 228954 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 229574 707718
rect 228954 707398 229574 707482
rect 228954 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 229574 707398
rect 228954 698614 229574 707162
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 266614 229574 302058
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 230614 229574 266058
rect 232674 708678 233294 711590
rect 232674 708442 232706 708678
rect 232942 708442 233026 708678
rect 233262 708442 233294 708678
rect 232674 708358 233294 708442
rect 232674 708122 232706 708358
rect 232942 708122 233026 708358
rect 233262 708122 233294 708358
rect 232674 666334 233294 708122
rect 232674 666098 232706 666334
rect 232942 666098 233026 666334
rect 233262 666098 233294 666334
rect 232674 666014 233294 666098
rect 232674 665778 232706 666014
rect 232942 665778 233026 666014
rect 233262 665778 233294 666014
rect 232674 630334 233294 665778
rect 232674 630098 232706 630334
rect 232942 630098 233026 630334
rect 233262 630098 233294 630334
rect 232674 630014 233294 630098
rect 232674 629778 232706 630014
rect 232942 629778 233026 630014
rect 233262 629778 233294 630014
rect 232674 594334 233294 629778
rect 232674 594098 232706 594334
rect 232942 594098 233026 594334
rect 233262 594098 233294 594334
rect 232674 594014 233294 594098
rect 232674 593778 232706 594014
rect 232942 593778 233026 594014
rect 233262 593778 233294 594014
rect 232674 558334 233294 593778
rect 232674 558098 232706 558334
rect 232942 558098 233026 558334
rect 233262 558098 233294 558334
rect 232674 558014 233294 558098
rect 232674 557778 232706 558014
rect 232942 557778 233026 558014
rect 233262 557778 233294 558014
rect 232674 522334 233294 557778
rect 232674 522098 232706 522334
rect 232942 522098 233026 522334
rect 233262 522098 233294 522334
rect 232674 522014 233294 522098
rect 232674 521778 232706 522014
rect 232942 521778 233026 522014
rect 233262 521778 233294 522014
rect 232674 486334 233294 521778
rect 232674 486098 232706 486334
rect 232942 486098 233026 486334
rect 233262 486098 233294 486334
rect 232674 486014 233294 486098
rect 232674 485778 232706 486014
rect 232942 485778 233026 486014
rect 233262 485778 233294 486014
rect 232674 450334 233294 485778
rect 232674 450098 232706 450334
rect 232942 450098 233026 450334
rect 233262 450098 233294 450334
rect 232674 450014 233294 450098
rect 232674 449778 232706 450014
rect 232942 449778 233026 450014
rect 233262 449778 233294 450014
rect 232674 414334 233294 449778
rect 232674 414098 232706 414334
rect 232942 414098 233026 414334
rect 233262 414098 233294 414334
rect 232674 414014 233294 414098
rect 232674 413778 232706 414014
rect 232942 413778 233026 414014
rect 233262 413778 233294 414014
rect 232674 378334 233294 413778
rect 232674 378098 232706 378334
rect 232942 378098 233026 378334
rect 233262 378098 233294 378334
rect 232674 378014 233294 378098
rect 232674 377778 232706 378014
rect 232942 377778 233026 378014
rect 233262 377778 233294 378014
rect 232674 342334 233294 377778
rect 232674 342098 232706 342334
rect 232942 342098 233026 342334
rect 233262 342098 233294 342334
rect 232674 342014 233294 342098
rect 232674 341778 232706 342014
rect 232942 341778 233026 342014
rect 233262 341778 233294 342014
rect 232674 306334 233294 341778
rect 232674 306098 232706 306334
rect 232942 306098 233026 306334
rect 233262 306098 233294 306334
rect 232674 306014 233294 306098
rect 232674 305778 232706 306014
rect 232942 305778 233026 306014
rect 233262 305778 233294 306014
rect 232674 270334 233294 305778
rect 232674 270098 232706 270334
rect 232942 270098 233026 270334
rect 233262 270098 233294 270334
rect 232674 270014 233294 270098
rect 232674 269778 232706 270014
rect 232942 269778 233026 270014
rect 233262 269778 233294 270014
rect 230427 240276 230493 240277
rect 230427 240212 230428 240276
rect 230492 240212 230493 240276
rect 230427 240211 230493 240212
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 230430 217973 230490 240211
rect 232674 234334 233294 269778
rect 232674 234098 232706 234334
rect 232942 234098 233026 234334
rect 233262 234098 233294 234334
rect 232674 234014 233294 234098
rect 232674 233778 232706 234014
rect 232942 233778 233026 234014
rect 233262 233778 233294 234014
rect 231899 227764 231965 227765
rect 231899 227700 231900 227764
rect 231964 227700 231965 227764
rect 231899 227699 231965 227700
rect 230427 217972 230493 217973
rect 230427 217908 230428 217972
rect 230492 217908 230493 217972
rect 230427 217907 230493 217908
rect 231902 204781 231962 227699
rect 231899 204780 231965 204781
rect 231899 204716 231900 204780
rect 231964 204716 231965 204780
rect 231899 204715 231965 204716
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 158614 229574 194058
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 228954 -3226 229574 14058
rect 228954 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 229574 -3226
rect 228954 -3546 229574 -3462
rect 228954 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 229574 -3546
rect 228954 -7654 229574 -3782
rect 232674 198334 233294 233778
rect 232674 198098 232706 198334
rect 232942 198098 233026 198334
rect 233262 198098 233294 198334
rect 232674 198014 233294 198098
rect 232674 197778 232706 198014
rect 232942 197778 233026 198014
rect 233262 197778 233294 198014
rect 232674 162334 233294 197778
rect 232674 162098 232706 162334
rect 232942 162098 233026 162334
rect 233262 162098 233294 162334
rect 232674 162014 233294 162098
rect 232674 161778 232706 162014
rect 232942 161778 233026 162014
rect 233262 161778 233294 162014
rect 232674 126334 233294 161778
rect 232674 126098 232706 126334
rect 232942 126098 233026 126334
rect 233262 126098 233294 126334
rect 232674 126014 233294 126098
rect 232674 125778 232706 126014
rect 232942 125778 233026 126014
rect 233262 125778 233294 126014
rect 232674 90334 233294 125778
rect 232674 90098 232706 90334
rect 232942 90098 233026 90334
rect 233262 90098 233294 90334
rect 232674 90014 233294 90098
rect 232674 89778 232706 90014
rect 232942 89778 233026 90014
rect 233262 89778 233294 90014
rect 232674 54334 233294 89778
rect 232674 54098 232706 54334
rect 232942 54098 233026 54334
rect 233262 54098 233294 54334
rect 232674 54014 233294 54098
rect 232674 53778 232706 54014
rect 232942 53778 233026 54014
rect 233262 53778 233294 54014
rect 232674 18334 233294 53778
rect 232674 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 233294 18334
rect 232674 18014 233294 18098
rect 232674 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 233294 18014
rect 232674 -4186 233294 17778
rect 232674 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 233294 -4186
rect 232674 -4506 233294 -4422
rect 232674 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 233294 -4506
rect 232674 -7654 233294 -4742
rect 236394 709638 237014 711590
rect 236394 709402 236426 709638
rect 236662 709402 236746 709638
rect 236982 709402 237014 709638
rect 236394 709318 237014 709402
rect 236394 709082 236426 709318
rect 236662 709082 236746 709318
rect 236982 709082 237014 709318
rect 236394 670054 237014 709082
rect 236394 669818 236426 670054
rect 236662 669818 236746 670054
rect 236982 669818 237014 670054
rect 236394 669734 237014 669818
rect 236394 669498 236426 669734
rect 236662 669498 236746 669734
rect 236982 669498 237014 669734
rect 236394 634054 237014 669498
rect 236394 633818 236426 634054
rect 236662 633818 236746 634054
rect 236982 633818 237014 634054
rect 236394 633734 237014 633818
rect 236394 633498 236426 633734
rect 236662 633498 236746 633734
rect 236982 633498 237014 633734
rect 236394 598054 237014 633498
rect 236394 597818 236426 598054
rect 236662 597818 236746 598054
rect 236982 597818 237014 598054
rect 236394 597734 237014 597818
rect 236394 597498 236426 597734
rect 236662 597498 236746 597734
rect 236982 597498 237014 597734
rect 236394 562054 237014 597498
rect 236394 561818 236426 562054
rect 236662 561818 236746 562054
rect 236982 561818 237014 562054
rect 236394 561734 237014 561818
rect 236394 561498 236426 561734
rect 236662 561498 236746 561734
rect 236982 561498 237014 561734
rect 236394 526054 237014 561498
rect 236394 525818 236426 526054
rect 236662 525818 236746 526054
rect 236982 525818 237014 526054
rect 236394 525734 237014 525818
rect 236394 525498 236426 525734
rect 236662 525498 236746 525734
rect 236982 525498 237014 525734
rect 236394 490054 237014 525498
rect 236394 489818 236426 490054
rect 236662 489818 236746 490054
rect 236982 489818 237014 490054
rect 236394 489734 237014 489818
rect 236394 489498 236426 489734
rect 236662 489498 236746 489734
rect 236982 489498 237014 489734
rect 236394 454054 237014 489498
rect 236394 453818 236426 454054
rect 236662 453818 236746 454054
rect 236982 453818 237014 454054
rect 236394 453734 237014 453818
rect 236394 453498 236426 453734
rect 236662 453498 236746 453734
rect 236982 453498 237014 453734
rect 236394 418054 237014 453498
rect 236394 417818 236426 418054
rect 236662 417818 236746 418054
rect 236982 417818 237014 418054
rect 236394 417734 237014 417818
rect 236394 417498 236426 417734
rect 236662 417498 236746 417734
rect 236982 417498 237014 417734
rect 236394 382054 237014 417498
rect 236394 381818 236426 382054
rect 236662 381818 236746 382054
rect 236982 381818 237014 382054
rect 236394 381734 237014 381818
rect 236394 381498 236426 381734
rect 236662 381498 236746 381734
rect 236982 381498 237014 381734
rect 236394 346054 237014 381498
rect 236394 345818 236426 346054
rect 236662 345818 236746 346054
rect 236982 345818 237014 346054
rect 236394 345734 237014 345818
rect 236394 345498 236426 345734
rect 236662 345498 236746 345734
rect 236982 345498 237014 345734
rect 236394 310054 237014 345498
rect 236394 309818 236426 310054
rect 236662 309818 236746 310054
rect 236982 309818 237014 310054
rect 236394 309734 237014 309818
rect 236394 309498 236426 309734
rect 236662 309498 236746 309734
rect 236982 309498 237014 309734
rect 236394 274054 237014 309498
rect 236394 273818 236426 274054
rect 236662 273818 236746 274054
rect 236982 273818 237014 274054
rect 236394 273734 237014 273818
rect 236394 273498 236426 273734
rect 236662 273498 236746 273734
rect 236982 273498 237014 273734
rect 236394 238054 237014 273498
rect 236394 237818 236426 238054
rect 236662 237818 236746 238054
rect 236982 237818 237014 238054
rect 236394 237734 237014 237818
rect 236394 237498 236426 237734
rect 236662 237498 236746 237734
rect 236982 237498 237014 237734
rect 236394 202054 237014 237498
rect 236394 201818 236426 202054
rect 236662 201818 236746 202054
rect 236982 201818 237014 202054
rect 236394 201734 237014 201818
rect 236394 201498 236426 201734
rect 236662 201498 236746 201734
rect 236982 201498 237014 201734
rect 236394 166054 237014 201498
rect 236394 165818 236426 166054
rect 236662 165818 236746 166054
rect 236982 165818 237014 166054
rect 236394 165734 237014 165818
rect 236394 165498 236426 165734
rect 236662 165498 236746 165734
rect 236982 165498 237014 165734
rect 236394 130054 237014 165498
rect 236394 129818 236426 130054
rect 236662 129818 236746 130054
rect 236982 129818 237014 130054
rect 236394 129734 237014 129818
rect 236394 129498 236426 129734
rect 236662 129498 236746 129734
rect 236982 129498 237014 129734
rect 236394 94054 237014 129498
rect 236394 93818 236426 94054
rect 236662 93818 236746 94054
rect 236982 93818 237014 94054
rect 236394 93734 237014 93818
rect 236394 93498 236426 93734
rect 236662 93498 236746 93734
rect 236982 93498 237014 93734
rect 236394 58054 237014 93498
rect 236394 57818 236426 58054
rect 236662 57818 236746 58054
rect 236982 57818 237014 58054
rect 236394 57734 237014 57818
rect 236394 57498 236426 57734
rect 236662 57498 236746 57734
rect 236982 57498 237014 57734
rect 236394 22054 237014 57498
rect 236394 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 237014 22054
rect 236394 21734 237014 21818
rect 236394 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 237014 21734
rect 236394 -5146 237014 21498
rect 236394 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 237014 -5146
rect 236394 -5466 237014 -5382
rect 236394 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 237014 -5466
rect 236394 -7654 237014 -5702
rect 240114 710598 240734 711590
rect 240114 710362 240146 710598
rect 240382 710362 240466 710598
rect 240702 710362 240734 710598
rect 240114 710278 240734 710362
rect 240114 710042 240146 710278
rect 240382 710042 240466 710278
rect 240702 710042 240734 710278
rect 240114 673774 240734 710042
rect 240114 673538 240146 673774
rect 240382 673538 240466 673774
rect 240702 673538 240734 673774
rect 240114 673454 240734 673538
rect 240114 673218 240146 673454
rect 240382 673218 240466 673454
rect 240702 673218 240734 673454
rect 240114 637774 240734 673218
rect 240114 637538 240146 637774
rect 240382 637538 240466 637774
rect 240702 637538 240734 637774
rect 240114 637454 240734 637538
rect 240114 637218 240146 637454
rect 240382 637218 240466 637454
rect 240702 637218 240734 637454
rect 240114 601774 240734 637218
rect 240114 601538 240146 601774
rect 240382 601538 240466 601774
rect 240702 601538 240734 601774
rect 240114 601454 240734 601538
rect 240114 601218 240146 601454
rect 240382 601218 240466 601454
rect 240702 601218 240734 601454
rect 240114 565774 240734 601218
rect 240114 565538 240146 565774
rect 240382 565538 240466 565774
rect 240702 565538 240734 565774
rect 240114 565454 240734 565538
rect 240114 565218 240146 565454
rect 240382 565218 240466 565454
rect 240702 565218 240734 565454
rect 240114 529774 240734 565218
rect 240114 529538 240146 529774
rect 240382 529538 240466 529774
rect 240702 529538 240734 529774
rect 240114 529454 240734 529538
rect 240114 529218 240146 529454
rect 240382 529218 240466 529454
rect 240702 529218 240734 529454
rect 240114 493774 240734 529218
rect 240114 493538 240146 493774
rect 240382 493538 240466 493774
rect 240702 493538 240734 493774
rect 240114 493454 240734 493538
rect 240114 493218 240146 493454
rect 240382 493218 240466 493454
rect 240702 493218 240734 493454
rect 240114 457774 240734 493218
rect 240114 457538 240146 457774
rect 240382 457538 240466 457774
rect 240702 457538 240734 457774
rect 240114 457454 240734 457538
rect 240114 457218 240146 457454
rect 240382 457218 240466 457454
rect 240702 457218 240734 457454
rect 240114 421774 240734 457218
rect 240114 421538 240146 421774
rect 240382 421538 240466 421774
rect 240702 421538 240734 421774
rect 240114 421454 240734 421538
rect 240114 421218 240146 421454
rect 240382 421218 240466 421454
rect 240702 421218 240734 421454
rect 240114 385774 240734 421218
rect 240114 385538 240146 385774
rect 240382 385538 240466 385774
rect 240702 385538 240734 385774
rect 240114 385454 240734 385538
rect 240114 385218 240146 385454
rect 240382 385218 240466 385454
rect 240702 385218 240734 385454
rect 240114 349774 240734 385218
rect 240114 349538 240146 349774
rect 240382 349538 240466 349774
rect 240702 349538 240734 349774
rect 240114 349454 240734 349538
rect 240114 349218 240146 349454
rect 240382 349218 240466 349454
rect 240702 349218 240734 349454
rect 240114 313774 240734 349218
rect 240114 313538 240146 313774
rect 240382 313538 240466 313774
rect 240702 313538 240734 313774
rect 240114 313454 240734 313538
rect 240114 313218 240146 313454
rect 240382 313218 240466 313454
rect 240702 313218 240734 313454
rect 240114 277774 240734 313218
rect 240114 277538 240146 277774
rect 240382 277538 240466 277774
rect 240702 277538 240734 277774
rect 240114 277454 240734 277538
rect 240114 277218 240146 277454
rect 240382 277218 240466 277454
rect 240702 277218 240734 277454
rect 240114 241774 240734 277218
rect 240114 241538 240146 241774
rect 240382 241538 240466 241774
rect 240702 241538 240734 241774
rect 240114 241454 240734 241538
rect 240114 241218 240146 241454
rect 240382 241218 240466 241454
rect 240702 241218 240734 241454
rect 240114 205774 240734 241218
rect 240114 205538 240146 205774
rect 240382 205538 240466 205774
rect 240702 205538 240734 205774
rect 240114 205454 240734 205538
rect 240114 205218 240146 205454
rect 240382 205218 240466 205454
rect 240702 205218 240734 205454
rect 240114 169774 240734 205218
rect 240114 169538 240146 169774
rect 240382 169538 240466 169774
rect 240702 169538 240734 169774
rect 240114 169454 240734 169538
rect 240114 169218 240146 169454
rect 240382 169218 240466 169454
rect 240702 169218 240734 169454
rect 240114 133774 240734 169218
rect 240114 133538 240146 133774
rect 240382 133538 240466 133774
rect 240702 133538 240734 133774
rect 240114 133454 240734 133538
rect 240114 133218 240146 133454
rect 240382 133218 240466 133454
rect 240702 133218 240734 133454
rect 240114 97774 240734 133218
rect 240114 97538 240146 97774
rect 240382 97538 240466 97774
rect 240702 97538 240734 97774
rect 240114 97454 240734 97538
rect 240114 97218 240146 97454
rect 240382 97218 240466 97454
rect 240702 97218 240734 97454
rect 240114 61774 240734 97218
rect 240114 61538 240146 61774
rect 240382 61538 240466 61774
rect 240702 61538 240734 61774
rect 240114 61454 240734 61538
rect 240114 61218 240146 61454
rect 240382 61218 240466 61454
rect 240702 61218 240734 61454
rect 240114 25774 240734 61218
rect 240114 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 240734 25774
rect 240114 25454 240734 25538
rect 240114 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 240734 25454
rect 240114 -6106 240734 25218
rect 240114 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 240734 -6106
rect 240114 -6426 240734 -6342
rect 240114 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 240734 -6426
rect 240114 -7654 240734 -6662
rect 243834 711558 244454 711590
rect 243834 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 244454 711558
rect 243834 711238 244454 711322
rect 243834 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 244454 711238
rect 243834 677494 244454 711002
rect 243834 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 244454 677494
rect 243834 677174 244454 677258
rect 243834 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 244454 677174
rect 243834 641494 244454 676938
rect 243834 641258 243866 641494
rect 244102 641258 244186 641494
rect 244422 641258 244454 641494
rect 243834 641174 244454 641258
rect 243834 640938 243866 641174
rect 244102 640938 244186 641174
rect 244422 640938 244454 641174
rect 243834 605494 244454 640938
rect 243834 605258 243866 605494
rect 244102 605258 244186 605494
rect 244422 605258 244454 605494
rect 243834 605174 244454 605258
rect 243834 604938 243866 605174
rect 244102 604938 244186 605174
rect 244422 604938 244454 605174
rect 243834 569494 244454 604938
rect 243834 569258 243866 569494
rect 244102 569258 244186 569494
rect 244422 569258 244454 569494
rect 243834 569174 244454 569258
rect 243834 568938 243866 569174
rect 244102 568938 244186 569174
rect 244422 568938 244454 569174
rect 243834 533494 244454 568938
rect 243834 533258 243866 533494
rect 244102 533258 244186 533494
rect 244422 533258 244454 533494
rect 243834 533174 244454 533258
rect 243834 532938 243866 533174
rect 244102 532938 244186 533174
rect 244422 532938 244454 533174
rect 243834 497494 244454 532938
rect 243834 497258 243866 497494
rect 244102 497258 244186 497494
rect 244422 497258 244454 497494
rect 243834 497174 244454 497258
rect 243834 496938 243866 497174
rect 244102 496938 244186 497174
rect 244422 496938 244454 497174
rect 243834 461494 244454 496938
rect 243834 461258 243866 461494
rect 244102 461258 244186 461494
rect 244422 461258 244454 461494
rect 243834 461174 244454 461258
rect 243834 460938 243866 461174
rect 244102 460938 244186 461174
rect 244422 460938 244454 461174
rect 243834 425494 244454 460938
rect 243834 425258 243866 425494
rect 244102 425258 244186 425494
rect 244422 425258 244454 425494
rect 243834 425174 244454 425258
rect 243834 424938 243866 425174
rect 244102 424938 244186 425174
rect 244422 424938 244454 425174
rect 243834 389494 244454 424938
rect 243834 389258 243866 389494
rect 244102 389258 244186 389494
rect 244422 389258 244454 389494
rect 243834 389174 244454 389258
rect 243834 388938 243866 389174
rect 244102 388938 244186 389174
rect 244422 388938 244454 389174
rect 243834 353494 244454 388938
rect 243834 353258 243866 353494
rect 244102 353258 244186 353494
rect 244422 353258 244454 353494
rect 243834 353174 244454 353258
rect 243834 352938 243866 353174
rect 244102 352938 244186 353174
rect 244422 352938 244454 353174
rect 243834 317494 244454 352938
rect 243834 317258 243866 317494
rect 244102 317258 244186 317494
rect 244422 317258 244454 317494
rect 243834 317174 244454 317258
rect 243834 316938 243866 317174
rect 244102 316938 244186 317174
rect 244422 316938 244454 317174
rect 243834 281494 244454 316938
rect 243834 281258 243866 281494
rect 244102 281258 244186 281494
rect 244422 281258 244454 281494
rect 243834 281174 244454 281258
rect 243834 280938 243866 281174
rect 244102 280938 244186 281174
rect 244422 280938 244454 281174
rect 243834 245494 244454 280938
rect 243834 245258 243866 245494
rect 244102 245258 244186 245494
rect 244422 245258 244454 245494
rect 243834 245174 244454 245258
rect 243834 244938 243866 245174
rect 244102 244938 244186 245174
rect 244422 244938 244454 245174
rect 243834 209494 244454 244938
rect 243834 209258 243866 209494
rect 244102 209258 244186 209494
rect 244422 209258 244454 209494
rect 243834 209174 244454 209258
rect 243834 208938 243866 209174
rect 244102 208938 244186 209174
rect 244422 208938 244454 209174
rect 243834 173494 244454 208938
rect 243834 173258 243866 173494
rect 244102 173258 244186 173494
rect 244422 173258 244454 173494
rect 243834 173174 244454 173258
rect 243834 172938 243866 173174
rect 244102 172938 244186 173174
rect 244422 172938 244454 173174
rect 243834 137494 244454 172938
rect 243834 137258 243866 137494
rect 244102 137258 244186 137494
rect 244422 137258 244454 137494
rect 243834 137174 244454 137258
rect 243834 136938 243866 137174
rect 244102 136938 244186 137174
rect 244422 136938 244454 137174
rect 243834 101494 244454 136938
rect 243834 101258 243866 101494
rect 244102 101258 244186 101494
rect 244422 101258 244454 101494
rect 243834 101174 244454 101258
rect 243834 100938 243866 101174
rect 244102 100938 244186 101174
rect 244422 100938 244454 101174
rect 243834 65494 244454 100938
rect 243834 65258 243866 65494
rect 244102 65258 244186 65494
rect 244422 65258 244454 65494
rect 243834 65174 244454 65258
rect 243834 64938 243866 65174
rect 244102 64938 244186 65174
rect 244422 64938 244454 65174
rect 243834 29494 244454 64938
rect 243834 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 244454 29494
rect 243834 29174 244454 29258
rect 243834 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 244454 29174
rect 243834 -7066 244454 28938
rect 243834 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 244454 -7066
rect 243834 -7386 244454 -7302
rect 243834 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 244454 -7386
rect 243834 -7654 244454 -7622
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 257514 705798 258134 711590
rect 257514 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 258134 705798
rect 257514 705478 258134 705562
rect 257514 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 258134 705478
rect 257514 691174 258134 705242
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 295174 258134 330618
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -1306 258134 6618
rect 257514 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 258134 -1306
rect 257514 -1626 258134 -1542
rect 257514 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 258134 -1626
rect 257514 -7654 258134 -1862
rect 261234 706758 261854 711590
rect 261234 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 261854 706758
rect 261234 706438 261854 706522
rect 261234 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 261854 706438
rect 261234 694894 261854 706202
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -2266 261854 10338
rect 261234 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 261854 -2266
rect 261234 -2586 261854 -2502
rect 261234 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 261854 -2586
rect 261234 -7654 261854 -2822
rect 264954 707718 265574 711590
rect 264954 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 265574 707718
rect 264954 707398 265574 707482
rect 264954 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 265574 707398
rect 264954 698614 265574 707162
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 264954 -3226 265574 14058
rect 264954 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 265574 -3226
rect 264954 -3546 265574 -3462
rect 264954 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 265574 -3546
rect 264954 -7654 265574 -3782
rect 268674 708678 269294 711590
rect 268674 708442 268706 708678
rect 268942 708442 269026 708678
rect 269262 708442 269294 708678
rect 268674 708358 269294 708442
rect 268674 708122 268706 708358
rect 268942 708122 269026 708358
rect 269262 708122 269294 708358
rect 268674 666334 269294 708122
rect 268674 666098 268706 666334
rect 268942 666098 269026 666334
rect 269262 666098 269294 666334
rect 268674 666014 269294 666098
rect 268674 665778 268706 666014
rect 268942 665778 269026 666014
rect 269262 665778 269294 666014
rect 268674 630334 269294 665778
rect 268674 630098 268706 630334
rect 268942 630098 269026 630334
rect 269262 630098 269294 630334
rect 268674 630014 269294 630098
rect 268674 629778 268706 630014
rect 268942 629778 269026 630014
rect 269262 629778 269294 630014
rect 268674 594334 269294 629778
rect 268674 594098 268706 594334
rect 268942 594098 269026 594334
rect 269262 594098 269294 594334
rect 268674 594014 269294 594098
rect 268674 593778 268706 594014
rect 268942 593778 269026 594014
rect 269262 593778 269294 594014
rect 268674 558334 269294 593778
rect 268674 558098 268706 558334
rect 268942 558098 269026 558334
rect 269262 558098 269294 558334
rect 268674 558014 269294 558098
rect 268674 557778 268706 558014
rect 268942 557778 269026 558014
rect 269262 557778 269294 558014
rect 268674 522334 269294 557778
rect 268674 522098 268706 522334
rect 268942 522098 269026 522334
rect 269262 522098 269294 522334
rect 268674 522014 269294 522098
rect 268674 521778 268706 522014
rect 268942 521778 269026 522014
rect 269262 521778 269294 522014
rect 268674 486334 269294 521778
rect 268674 486098 268706 486334
rect 268942 486098 269026 486334
rect 269262 486098 269294 486334
rect 268674 486014 269294 486098
rect 268674 485778 268706 486014
rect 268942 485778 269026 486014
rect 269262 485778 269294 486014
rect 268674 450334 269294 485778
rect 268674 450098 268706 450334
rect 268942 450098 269026 450334
rect 269262 450098 269294 450334
rect 268674 450014 269294 450098
rect 268674 449778 268706 450014
rect 268942 449778 269026 450014
rect 269262 449778 269294 450014
rect 268674 414334 269294 449778
rect 268674 414098 268706 414334
rect 268942 414098 269026 414334
rect 269262 414098 269294 414334
rect 268674 414014 269294 414098
rect 268674 413778 268706 414014
rect 268942 413778 269026 414014
rect 269262 413778 269294 414014
rect 268674 378334 269294 413778
rect 268674 378098 268706 378334
rect 268942 378098 269026 378334
rect 269262 378098 269294 378334
rect 268674 378014 269294 378098
rect 268674 377778 268706 378014
rect 268942 377778 269026 378014
rect 269262 377778 269294 378014
rect 268674 342334 269294 377778
rect 268674 342098 268706 342334
rect 268942 342098 269026 342334
rect 269262 342098 269294 342334
rect 268674 342014 269294 342098
rect 268674 341778 268706 342014
rect 268942 341778 269026 342014
rect 269262 341778 269294 342014
rect 268674 306334 269294 341778
rect 268674 306098 268706 306334
rect 268942 306098 269026 306334
rect 269262 306098 269294 306334
rect 268674 306014 269294 306098
rect 268674 305778 268706 306014
rect 268942 305778 269026 306014
rect 269262 305778 269294 306014
rect 268674 270334 269294 305778
rect 268674 270098 268706 270334
rect 268942 270098 269026 270334
rect 269262 270098 269294 270334
rect 268674 270014 269294 270098
rect 268674 269778 268706 270014
rect 268942 269778 269026 270014
rect 269262 269778 269294 270014
rect 268674 234334 269294 269778
rect 268674 234098 268706 234334
rect 268942 234098 269026 234334
rect 269262 234098 269294 234334
rect 268674 234014 269294 234098
rect 268674 233778 268706 234014
rect 268942 233778 269026 234014
rect 269262 233778 269294 234014
rect 268674 198334 269294 233778
rect 268674 198098 268706 198334
rect 268942 198098 269026 198334
rect 269262 198098 269294 198334
rect 268674 198014 269294 198098
rect 268674 197778 268706 198014
rect 268942 197778 269026 198014
rect 269262 197778 269294 198014
rect 268674 162334 269294 197778
rect 268674 162098 268706 162334
rect 268942 162098 269026 162334
rect 269262 162098 269294 162334
rect 268674 162014 269294 162098
rect 268674 161778 268706 162014
rect 268942 161778 269026 162014
rect 269262 161778 269294 162014
rect 268674 126334 269294 161778
rect 268674 126098 268706 126334
rect 268942 126098 269026 126334
rect 269262 126098 269294 126334
rect 268674 126014 269294 126098
rect 268674 125778 268706 126014
rect 268942 125778 269026 126014
rect 269262 125778 269294 126014
rect 268674 90334 269294 125778
rect 268674 90098 268706 90334
rect 268942 90098 269026 90334
rect 269262 90098 269294 90334
rect 268674 90014 269294 90098
rect 268674 89778 268706 90014
rect 268942 89778 269026 90014
rect 269262 89778 269294 90014
rect 268674 54334 269294 89778
rect 268674 54098 268706 54334
rect 268942 54098 269026 54334
rect 269262 54098 269294 54334
rect 268674 54014 269294 54098
rect 268674 53778 268706 54014
rect 268942 53778 269026 54014
rect 269262 53778 269294 54014
rect 268674 18334 269294 53778
rect 268674 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 269294 18334
rect 268674 18014 269294 18098
rect 268674 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 269294 18014
rect 268674 -4186 269294 17778
rect 268674 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 269294 -4186
rect 268674 -4506 269294 -4422
rect 268674 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 269294 -4506
rect 268674 -7654 269294 -4742
rect 272394 709638 273014 711590
rect 272394 709402 272426 709638
rect 272662 709402 272746 709638
rect 272982 709402 273014 709638
rect 272394 709318 273014 709402
rect 272394 709082 272426 709318
rect 272662 709082 272746 709318
rect 272982 709082 273014 709318
rect 272394 670054 273014 709082
rect 272394 669818 272426 670054
rect 272662 669818 272746 670054
rect 272982 669818 273014 670054
rect 272394 669734 273014 669818
rect 272394 669498 272426 669734
rect 272662 669498 272746 669734
rect 272982 669498 273014 669734
rect 272394 634054 273014 669498
rect 272394 633818 272426 634054
rect 272662 633818 272746 634054
rect 272982 633818 273014 634054
rect 272394 633734 273014 633818
rect 272394 633498 272426 633734
rect 272662 633498 272746 633734
rect 272982 633498 273014 633734
rect 272394 598054 273014 633498
rect 272394 597818 272426 598054
rect 272662 597818 272746 598054
rect 272982 597818 273014 598054
rect 272394 597734 273014 597818
rect 272394 597498 272426 597734
rect 272662 597498 272746 597734
rect 272982 597498 273014 597734
rect 272394 562054 273014 597498
rect 272394 561818 272426 562054
rect 272662 561818 272746 562054
rect 272982 561818 273014 562054
rect 272394 561734 273014 561818
rect 272394 561498 272426 561734
rect 272662 561498 272746 561734
rect 272982 561498 273014 561734
rect 272394 526054 273014 561498
rect 272394 525818 272426 526054
rect 272662 525818 272746 526054
rect 272982 525818 273014 526054
rect 272394 525734 273014 525818
rect 272394 525498 272426 525734
rect 272662 525498 272746 525734
rect 272982 525498 273014 525734
rect 272394 490054 273014 525498
rect 272394 489818 272426 490054
rect 272662 489818 272746 490054
rect 272982 489818 273014 490054
rect 272394 489734 273014 489818
rect 272394 489498 272426 489734
rect 272662 489498 272746 489734
rect 272982 489498 273014 489734
rect 272394 454054 273014 489498
rect 272394 453818 272426 454054
rect 272662 453818 272746 454054
rect 272982 453818 273014 454054
rect 272394 453734 273014 453818
rect 272394 453498 272426 453734
rect 272662 453498 272746 453734
rect 272982 453498 273014 453734
rect 272394 418054 273014 453498
rect 272394 417818 272426 418054
rect 272662 417818 272746 418054
rect 272982 417818 273014 418054
rect 272394 417734 273014 417818
rect 272394 417498 272426 417734
rect 272662 417498 272746 417734
rect 272982 417498 273014 417734
rect 272394 382054 273014 417498
rect 272394 381818 272426 382054
rect 272662 381818 272746 382054
rect 272982 381818 273014 382054
rect 272394 381734 273014 381818
rect 272394 381498 272426 381734
rect 272662 381498 272746 381734
rect 272982 381498 273014 381734
rect 272394 346054 273014 381498
rect 272394 345818 272426 346054
rect 272662 345818 272746 346054
rect 272982 345818 273014 346054
rect 272394 345734 273014 345818
rect 272394 345498 272426 345734
rect 272662 345498 272746 345734
rect 272982 345498 273014 345734
rect 272394 310054 273014 345498
rect 272394 309818 272426 310054
rect 272662 309818 272746 310054
rect 272982 309818 273014 310054
rect 272394 309734 273014 309818
rect 272394 309498 272426 309734
rect 272662 309498 272746 309734
rect 272982 309498 273014 309734
rect 272394 274054 273014 309498
rect 272394 273818 272426 274054
rect 272662 273818 272746 274054
rect 272982 273818 273014 274054
rect 272394 273734 273014 273818
rect 272394 273498 272426 273734
rect 272662 273498 272746 273734
rect 272982 273498 273014 273734
rect 272394 238054 273014 273498
rect 272394 237818 272426 238054
rect 272662 237818 272746 238054
rect 272982 237818 273014 238054
rect 272394 237734 273014 237818
rect 272394 237498 272426 237734
rect 272662 237498 272746 237734
rect 272982 237498 273014 237734
rect 272394 202054 273014 237498
rect 272394 201818 272426 202054
rect 272662 201818 272746 202054
rect 272982 201818 273014 202054
rect 272394 201734 273014 201818
rect 272394 201498 272426 201734
rect 272662 201498 272746 201734
rect 272982 201498 273014 201734
rect 272394 166054 273014 201498
rect 272394 165818 272426 166054
rect 272662 165818 272746 166054
rect 272982 165818 273014 166054
rect 272394 165734 273014 165818
rect 272394 165498 272426 165734
rect 272662 165498 272746 165734
rect 272982 165498 273014 165734
rect 272394 130054 273014 165498
rect 272394 129818 272426 130054
rect 272662 129818 272746 130054
rect 272982 129818 273014 130054
rect 272394 129734 273014 129818
rect 272394 129498 272426 129734
rect 272662 129498 272746 129734
rect 272982 129498 273014 129734
rect 272394 94054 273014 129498
rect 272394 93818 272426 94054
rect 272662 93818 272746 94054
rect 272982 93818 273014 94054
rect 272394 93734 273014 93818
rect 272394 93498 272426 93734
rect 272662 93498 272746 93734
rect 272982 93498 273014 93734
rect 272394 58054 273014 93498
rect 272394 57818 272426 58054
rect 272662 57818 272746 58054
rect 272982 57818 273014 58054
rect 272394 57734 273014 57818
rect 272394 57498 272426 57734
rect 272662 57498 272746 57734
rect 272982 57498 273014 57734
rect 272394 22054 273014 57498
rect 272394 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 273014 22054
rect 272394 21734 273014 21818
rect 272394 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 273014 21734
rect 272394 -5146 273014 21498
rect 272394 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 273014 -5146
rect 272394 -5466 273014 -5382
rect 272394 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 273014 -5466
rect 272394 -7654 273014 -5702
rect 276114 710598 276734 711590
rect 276114 710362 276146 710598
rect 276382 710362 276466 710598
rect 276702 710362 276734 710598
rect 276114 710278 276734 710362
rect 276114 710042 276146 710278
rect 276382 710042 276466 710278
rect 276702 710042 276734 710278
rect 276114 673774 276734 710042
rect 276114 673538 276146 673774
rect 276382 673538 276466 673774
rect 276702 673538 276734 673774
rect 276114 673454 276734 673538
rect 276114 673218 276146 673454
rect 276382 673218 276466 673454
rect 276702 673218 276734 673454
rect 276114 637774 276734 673218
rect 276114 637538 276146 637774
rect 276382 637538 276466 637774
rect 276702 637538 276734 637774
rect 276114 637454 276734 637538
rect 276114 637218 276146 637454
rect 276382 637218 276466 637454
rect 276702 637218 276734 637454
rect 276114 601774 276734 637218
rect 276114 601538 276146 601774
rect 276382 601538 276466 601774
rect 276702 601538 276734 601774
rect 276114 601454 276734 601538
rect 276114 601218 276146 601454
rect 276382 601218 276466 601454
rect 276702 601218 276734 601454
rect 276114 565774 276734 601218
rect 276114 565538 276146 565774
rect 276382 565538 276466 565774
rect 276702 565538 276734 565774
rect 276114 565454 276734 565538
rect 276114 565218 276146 565454
rect 276382 565218 276466 565454
rect 276702 565218 276734 565454
rect 276114 529774 276734 565218
rect 276114 529538 276146 529774
rect 276382 529538 276466 529774
rect 276702 529538 276734 529774
rect 276114 529454 276734 529538
rect 276114 529218 276146 529454
rect 276382 529218 276466 529454
rect 276702 529218 276734 529454
rect 276114 493774 276734 529218
rect 276114 493538 276146 493774
rect 276382 493538 276466 493774
rect 276702 493538 276734 493774
rect 276114 493454 276734 493538
rect 276114 493218 276146 493454
rect 276382 493218 276466 493454
rect 276702 493218 276734 493454
rect 276114 457774 276734 493218
rect 276114 457538 276146 457774
rect 276382 457538 276466 457774
rect 276702 457538 276734 457774
rect 276114 457454 276734 457538
rect 276114 457218 276146 457454
rect 276382 457218 276466 457454
rect 276702 457218 276734 457454
rect 276114 421774 276734 457218
rect 276114 421538 276146 421774
rect 276382 421538 276466 421774
rect 276702 421538 276734 421774
rect 276114 421454 276734 421538
rect 276114 421218 276146 421454
rect 276382 421218 276466 421454
rect 276702 421218 276734 421454
rect 276114 385774 276734 421218
rect 276114 385538 276146 385774
rect 276382 385538 276466 385774
rect 276702 385538 276734 385774
rect 276114 385454 276734 385538
rect 276114 385218 276146 385454
rect 276382 385218 276466 385454
rect 276702 385218 276734 385454
rect 276114 349774 276734 385218
rect 276114 349538 276146 349774
rect 276382 349538 276466 349774
rect 276702 349538 276734 349774
rect 276114 349454 276734 349538
rect 276114 349218 276146 349454
rect 276382 349218 276466 349454
rect 276702 349218 276734 349454
rect 276114 313774 276734 349218
rect 276114 313538 276146 313774
rect 276382 313538 276466 313774
rect 276702 313538 276734 313774
rect 276114 313454 276734 313538
rect 276114 313218 276146 313454
rect 276382 313218 276466 313454
rect 276702 313218 276734 313454
rect 276114 277774 276734 313218
rect 276114 277538 276146 277774
rect 276382 277538 276466 277774
rect 276702 277538 276734 277774
rect 276114 277454 276734 277538
rect 276114 277218 276146 277454
rect 276382 277218 276466 277454
rect 276702 277218 276734 277454
rect 276114 241774 276734 277218
rect 276114 241538 276146 241774
rect 276382 241538 276466 241774
rect 276702 241538 276734 241774
rect 276114 241454 276734 241538
rect 276114 241218 276146 241454
rect 276382 241218 276466 241454
rect 276702 241218 276734 241454
rect 276114 205774 276734 241218
rect 276114 205538 276146 205774
rect 276382 205538 276466 205774
rect 276702 205538 276734 205774
rect 276114 205454 276734 205538
rect 276114 205218 276146 205454
rect 276382 205218 276466 205454
rect 276702 205218 276734 205454
rect 276114 169774 276734 205218
rect 276114 169538 276146 169774
rect 276382 169538 276466 169774
rect 276702 169538 276734 169774
rect 276114 169454 276734 169538
rect 276114 169218 276146 169454
rect 276382 169218 276466 169454
rect 276702 169218 276734 169454
rect 276114 133774 276734 169218
rect 276114 133538 276146 133774
rect 276382 133538 276466 133774
rect 276702 133538 276734 133774
rect 276114 133454 276734 133538
rect 276114 133218 276146 133454
rect 276382 133218 276466 133454
rect 276702 133218 276734 133454
rect 276114 97774 276734 133218
rect 276114 97538 276146 97774
rect 276382 97538 276466 97774
rect 276702 97538 276734 97774
rect 276114 97454 276734 97538
rect 276114 97218 276146 97454
rect 276382 97218 276466 97454
rect 276702 97218 276734 97454
rect 276114 61774 276734 97218
rect 276114 61538 276146 61774
rect 276382 61538 276466 61774
rect 276702 61538 276734 61774
rect 276114 61454 276734 61538
rect 276114 61218 276146 61454
rect 276382 61218 276466 61454
rect 276702 61218 276734 61454
rect 276114 25774 276734 61218
rect 276114 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 276734 25774
rect 276114 25454 276734 25538
rect 276114 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 276734 25454
rect 276114 -6106 276734 25218
rect 276114 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 276734 -6106
rect 276114 -6426 276734 -6342
rect 276114 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 276734 -6426
rect 276114 -7654 276734 -6662
rect 279834 711558 280454 711590
rect 279834 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 280454 711558
rect 279834 711238 280454 711322
rect 279834 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 280454 711238
rect 279834 677494 280454 711002
rect 279834 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 280454 677494
rect 279834 677174 280454 677258
rect 279834 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 280454 677174
rect 279834 641494 280454 676938
rect 279834 641258 279866 641494
rect 280102 641258 280186 641494
rect 280422 641258 280454 641494
rect 279834 641174 280454 641258
rect 279834 640938 279866 641174
rect 280102 640938 280186 641174
rect 280422 640938 280454 641174
rect 279834 605494 280454 640938
rect 279834 605258 279866 605494
rect 280102 605258 280186 605494
rect 280422 605258 280454 605494
rect 279834 605174 280454 605258
rect 279834 604938 279866 605174
rect 280102 604938 280186 605174
rect 280422 604938 280454 605174
rect 279834 569494 280454 604938
rect 279834 569258 279866 569494
rect 280102 569258 280186 569494
rect 280422 569258 280454 569494
rect 279834 569174 280454 569258
rect 279834 568938 279866 569174
rect 280102 568938 280186 569174
rect 280422 568938 280454 569174
rect 279834 533494 280454 568938
rect 279834 533258 279866 533494
rect 280102 533258 280186 533494
rect 280422 533258 280454 533494
rect 279834 533174 280454 533258
rect 279834 532938 279866 533174
rect 280102 532938 280186 533174
rect 280422 532938 280454 533174
rect 279834 497494 280454 532938
rect 279834 497258 279866 497494
rect 280102 497258 280186 497494
rect 280422 497258 280454 497494
rect 279834 497174 280454 497258
rect 279834 496938 279866 497174
rect 280102 496938 280186 497174
rect 280422 496938 280454 497174
rect 279834 461494 280454 496938
rect 279834 461258 279866 461494
rect 280102 461258 280186 461494
rect 280422 461258 280454 461494
rect 279834 461174 280454 461258
rect 279834 460938 279866 461174
rect 280102 460938 280186 461174
rect 280422 460938 280454 461174
rect 279834 425494 280454 460938
rect 279834 425258 279866 425494
rect 280102 425258 280186 425494
rect 280422 425258 280454 425494
rect 279834 425174 280454 425258
rect 279834 424938 279866 425174
rect 280102 424938 280186 425174
rect 280422 424938 280454 425174
rect 279834 389494 280454 424938
rect 279834 389258 279866 389494
rect 280102 389258 280186 389494
rect 280422 389258 280454 389494
rect 279834 389174 280454 389258
rect 279834 388938 279866 389174
rect 280102 388938 280186 389174
rect 280422 388938 280454 389174
rect 279834 353494 280454 388938
rect 279834 353258 279866 353494
rect 280102 353258 280186 353494
rect 280422 353258 280454 353494
rect 279834 353174 280454 353258
rect 279834 352938 279866 353174
rect 280102 352938 280186 353174
rect 280422 352938 280454 353174
rect 279834 317494 280454 352938
rect 279834 317258 279866 317494
rect 280102 317258 280186 317494
rect 280422 317258 280454 317494
rect 279834 317174 280454 317258
rect 279834 316938 279866 317174
rect 280102 316938 280186 317174
rect 280422 316938 280454 317174
rect 279834 281494 280454 316938
rect 279834 281258 279866 281494
rect 280102 281258 280186 281494
rect 280422 281258 280454 281494
rect 279834 281174 280454 281258
rect 279834 280938 279866 281174
rect 280102 280938 280186 281174
rect 280422 280938 280454 281174
rect 279834 245494 280454 280938
rect 279834 245258 279866 245494
rect 280102 245258 280186 245494
rect 280422 245258 280454 245494
rect 279834 245174 280454 245258
rect 279834 244938 279866 245174
rect 280102 244938 280186 245174
rect 280422 244938 280454 245174
rect 279834 209494 280454 244938
rect 279834 209258 279866 209494
rect 280102 209258 280186 209494
rect 280422 209258 280454 209494
rect 279834 209174 280454 209258
rect 279834 208938 279866 209174
rect 280102 208938 280186 209174
rect 280422 208938 280454 209174
rect 279834 173494 280454 208938
rect 279834 173258 279866 173494
rect 280102 173258 280186 173494
rect 280422 173258 280454 173494
rect 279834 173174 280454 173258
rect 279834 172938 279866 173174
rect 280102 172938 280186 173174
rect 280422 172938 280454 173174
rect 279834 137494 280454 172938
rect 279834 137258 279866 137494
rect 280102 137258 280186 137494
rect 280422 137258 280454 137494
rect 279834 137174 280454 137258
rect 279834 136938 279866 137174
rect 280102 136938 280186 137174
rect 280422 136938 280454 137174
rect 279834 101494 280454 136938
rect 279834 101258 279866 101494
rect 280102 101258 280186 101494
rect 280422 101258 280454 101494
rect 279834 101174 280454 101258
rect 279834 100938 279866 101174
rect 280102 100938 280186 101174
rect 280422 100938 280454 101174
rect 279834 65494 280454 100938
rect 279834 65258 279866 65494
rect 280102 65258 280186 65494
rect 280422 65258 280454 65494
rect 279834 65174 280454 65258
rect 279834 64938 279866 65174
rect 280102 64938 280186 65174
rect 280422 64938 280454 65174
rect 279834 29494 280454 64938
rect 279834 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 280454 29494
rect 279834 29174 280454 29258
rect 279834 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 280454 29174
rect 279834 -7066 280454 28938
rect 279834 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 280454 -7066
rect 279834 -7386 280454 -7302
rect 279834 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 280454 -7386
rect 279834 -7654 280454 -7622
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 293514 705798 294134 711590
rect 293514 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 294134 705798
rect 293514 705478 294134 705562
rect 293514 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 294134 705478
rect 293514 691174 294134 705242
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -1306 294134 6618
rect 293514 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 294134 -1306
rect 293514 -1626 294134 -1542
rect 293514 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 294134 -1626
rect 293514 -7654 294134 -1862
rect 297234 706758 297854 711590
rect 297234 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 297854 706758
rect 297234 706438 297854 706522
rect 297234 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 297854 706438
rect 297234 694894 297854 706202
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -2266 297854 10338
rect 297234 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 297854 -2266
rect 297234 -2586 297854 -2502
rect 297234 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 297854 -2586
rect 297234 -7654 297854 -2822
rect 300954 707718 301574 711590
rect 300954 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 301574 707718
rect 300954 707398 301574 707482
rect 300954 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 301574 707398
rect 300954 698614 301574 707162
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 300954 -3226 301574 14058
rect 300954 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 301574 -3226
rect 300954 -3546 301574 -3462
rect 300954 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 301574 -3546
rect 300954 -7654 301574 -3782
rect 304674 708678 305294 711590
rect 304674 708442 304706 708678
rect 304942 708442 305026 708678
rect 305262 708442 305294 708678
rect 304674 708358 305294 708442
rect 304674 708122 304706 708358
rect 304942 708122 305026 708358
rect 305262 708122 305294 708358
rect 304674 666334 305294 708122
rect 304674 666098 304706 666334
rect 304942 666098 305026 666334
rect 305262 666098 305294 666334
rect 304674 666014 305294 666098
rect 304674 665778 304706 666014
rect 304942 665778 305026 666014
rect 305262 665778 305294 666014
rect 304674 630334 305294 665778
rect 304674 630098 304706 630334
rect 304942 630098 305026 630334
rect 305262 630098 305294 630334
rect 304674 630014 305294 630098
rect 304674 629778 304706 630014
rect 304942 629778 305026 630014
rect 305262 629778 305294 630014
rect 304674 594334 305294 629778
rect 304674 594098 304706 594334
rect 304942 594098 305026 594334
rect 305262 594098 305294 594334
rect 304674 594014 305294 594098
rect 304674 593778 304706 594014
rect 304942 593778 305026 594014
rect 305262 593778 305294 594014
rect 304674 558334 305294 593778
rect 304674 558098 304706 558334
rect 304942 558098 305026 558334
rect 305262 558098 305294 558334
rect 304674 558014 305294 558098
rect 304674 557778 304706 558014
rect 304942 557778 305026 558014
rect 305262 557778 305294 558014
rect 304674 522334 305294 557778
rect 304674 522098 304706 522334
rect 304942 522098 305026 522334
rect 305262 522098 305294 522334
rect 304674 522014 305294 522098
rect 304674 521778 304706 522014
rect 304942 521778 305026 522014
rect 305262 521778 305294 522014
rect 304674 486334 305294 521778
rect 304674 486098 304706 486334
rect 304942 486098 305026 486334
rect 305262 486098 305294 486334
rect 304674 486014 305294 486098
rect 304674 485778 304706 486014
rect 304942 485778 305026 486014
rect 305262 485778 305294 486014
rect 304674 450334 305294 485778
rect 304674 450098 304706 450334
rect 304942 450098 305026 450334
rect 305262 450098 305294 450334
rect 304674 450014 305294 450098
rect 304674 449778 304706 450014
rect 304942 449778 305026 450014
rect 305262 449778 305294 450014
rect 304674 414334 305294 449778
rect 304674 414098 304706 414334
rect 304942 414098 305026 414334
rect 305262 414098 305294 414334
rect 304674 414014 305294 414098
rect 304674 413778 304706 414014
rect 304942 413778 305026 414014
rect 305262 413778 305294 414014
rect 304674 378334 305294 413778
rect 304674 378098 304706 378334
rect 304942 378098 305026 378334
rect 305262 378098 305294 378334
rect 304674 378014 305294 378098
rect 304674 377778 304706 378014
rect 304942 377778 305026 378014
rect 305262 377778 305294 378014
rect 304674 342334 305294 377778
rect 304674 342098 304706 342334
rect 304942 342098 305026 342334
rect 305262 342098 305294 342334
rect 304674 342014 305294 342098
rect 304674 341778 304706 342014
rect 304942 341778 305026 342014
rect 305262 341778 305294 342014
rect 304674 306334 305294 341778
rect 304674 306098 304706 306334
rect 304942 306098 305026 306334
rect 305262 306098 305294 306334
rect 304674 306014 305294 306098
rect 304674 305778 304706 306014
rect 304942 305778 305026 306014
rect 305262 305778 305294 306014
rect 304674 270334 305294 305778
rect 304674 270098 304706 270334
rect 304942 270098 305026 270334
rect 305262 270098 305294 270334
rect 304674 270014 305294 270098
rect 304674 269778 304706 270014
rect 304942 269778 305026 270014
rect 305262 269778 305294 270014
rect 304674 234334 305294 269778
rect 304674 234098 304706 234334
rect 304942 234098 305026 234334
rect 305262 234098 305294 234334
rect 304674 234014 305294 234098
rect 304674 233778 304706 234014
rect 304942 233778 305026 234014
rect 305262 233778 305294 234014
rect 304674 198334 305294 233778
rect 304674 198098 304706 198334
rect 304942 198098 305026 198334
rect 305262 198098 305294 198334
rect 304674 198014 305294 198098
rect 304674 197778 304706 198014
rect 304942 197778 305026 198014
rect 305262 197778 305294 198014
rect 304674 162334 305294 197778
rect 304674 162098 304706 162334
rect 304942 162098 305026 162334
rect 305262 162098 305294 162334
rect 304674 162014 305294 162098
rect 304674 161778 304706 162014
rect 304942 161778 305026 162014
rect 305262 161778 305294 162014
rect 304674 126334 305294 161778
rect 304674 126098 304706 126334
rect 304942 126098 305026 126334
rect 305262 126098 305294 126334
rect 304674 126014 305294 126098
rect 304674 125778 304706 126014
rect 304942 125778 305026 126014
rect 305262 125778 305294 126014
rect 304674 90334 305294 125778
rect 304674 90098 304706 90334
rect 304942 90098 305026 90334
rect 305262 90098 305294 90334
rect 304674 90014 305294 90098
rect 304674 89778 304706 90014
rect 304942 89778 305026 90014
rect 305262 89778 305294 90014
rect 304674 54334 305294 89778
rect 304674 54098 304706 54334
rect 304942 54098 305026 54334
rect 305262 54098 305294 54334
rect 304674 54014 305294 54098
rect 304674 53778 304706 54014
rect 304942 53778 305026 54014
rect 305262 53778 305294 54014
rect 304674 18334 305294 53778
rect 304674 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 305294 18334
rect 304674 18014 305294 18098
rect 304674 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 305294 18014
rect 304674 -4186 305294 17778
rect 304674 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 305294 -4186
rect 304674 -4506 305294 -4422
rect 304674 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 305294 -4506
rect 304674 -7654 305294 -4742
rect 308394 709638 309014 711590
rect 308394 709402 308426 709638
rect 308662 709402 308746 709638
rect 308982 709402 309014 709638
rect 308394 709318 309014 709402
rect 308394 709082 308426 709318
rect 308662 709082 308746 709318
rect 308982 709082 309014 709318
rect 308394 670054 309014 709082
rect 308394 669818 308426 670054
rect 308662 669818 308746 670054
rect 308982 669818 309014 670054
rect 308394 669734 309014 669818
rect 308394 669498 308426 669734
rect 308662 669498 308746 669734
rect 308982 669498 309014 669734
rect 308394 634054 309014 669498
rect 308394 633818 308426 634054
rect 308662 633818 308746 634054
rect 308982 633818 309014 634054
rect 308394 633734 309014 633818
rect 308394 633498 308426 633734
rect 308662 633498 308746 633734
rect 308982 633498 309014 633734
rect 308394 598054 309014 633498
rect 308394 597818 308426 598054
rect 308662 597818 308746 598054
rect 308982 597818 309014 598054
rect 308394 597734 309014 597818
rect 308394 597498 308426 597734
rect 308662 597498 308746 597734
rect 308982 597498 309014 597734
rect 308394 562054 309014 597498
rect 308394 561818 308426 562054
rect 308662 561818 308746 562054
rect 308982 561818 309014 562054
rect 308394 561734 309014 561818
rect 308394 561498 308426 561734
rect 308662 561498 308746 561734
rect 308982 561498 309014 561734
rect 308394 526054 309014 561498
rect 308394 525818 308426 526054
rect 308662 525818 308746 526054
rect 308982 525818 309014 526054
rect 308394 525734 309014 525818
rect 308394 525498 308426 525734
rect 308662 525498 308746 525734
rect 308982 525498 309014 525734
rect 308394 490054 309014 525498
rect 308394 489818 308426 490054
rect 308662 489818 308746 490054
rect 308982 489818 309014 490054
rect 308394 489734 309014 489818
rect 308394 489498 308426 489734
rect 308662 489498 308746 489734
rect 308982 489498 309014 489734
rect 308394 454054 309014 489498
rect 308394 453818 308426 454054
rect 308662 453818 308746 454054
rect 308982 453818 309014 454054
rect 308394 453734 309014 453818
rect 308394 453498 308426 453734
rect 308662 453498 308746 453734
rect 308982 453498 309014 453734
rect 308394 418054 309014 453498
rect 308394 417818 308426 418054
rect 308662 417818 308746 418054
rect 308982 417818 309014 418054
rect 308394 417734 309014 417818
rect 308394 417498 308426 417734
rect 308662 417498 308746 417734
rect 308982 417498 309014 417734
rect 308394 382054 309014 417498
rect 308394 381818 308426 382054
rect 308662 381818 308746 382054
rect 308982 381818 309014 382054
rect 308394 381734 309014 381818
rect 308394 381498 308426 381734
rect 308662 381498 308746 381734
rect 308982 381498 309014 381734
rect 308394 346054 309014 381498
rect 308394 345818 308426 346054
rect 308662 345818 308746 346054
rect 308982 345818 309014 346054
rect 308394 345734 309014 345818
rect 308394 345498 308426 345734
rect 308662 345498 308746 345734
rect 308982 345498 309014 345734
rect 308394 310054 309014 345498
rect 308394 309818 308426 310054
rect 308662 309818 308746 310054
rect 308982 309818 309014 310054
rect 308394 309734 309014 309818
rect 308394 309498 308426 309734
rect 308662 309498 308746 309734
rect 308982 309498 309014 309734
rect 308394 274054 309014 309498
rect 308394 273818 308426 274054
rect 308662 273818 308746 274054
rect 308982 273818 309014 274054
rect 308394 273734 309014 273818
rect 308394 273498 308426 273734
rect 308662 273498 308746 273734
rect 308982 273498 309014 273734
rect 308394 238054 309014 273498
rect 308394 237818 308426 238054
rect 308662 237818 308746 238054
rect 308982 237818 309014 238054
rect 308394 237734 309014 237818
rect 308394 237498 308426 237734
rect 308662 237498 308746 237734
rect 308982 237498 309014 237734
rect 308394 202054 309014 237498
rect 308394 201818 308426 202054
rect 308662 201818 308746 202054
rect 308982 201818 309014 202054
rect 308394 201734 309014 201818
rect 308394 201498 308426 201734
rect 308662 201498 308746 201734
rect 308982 201498 309014 201734
rect 308394 166054 309014 201498
rect 308394 165818 308426 166054
rect 308662 165818 308746 166054
rect 308982 165818 309014 166054
rect 308394 165734 309014 165818
rect 308394 165498 308426 165734
rect 308662 165498 308746 165734
rect 308982 165498 309014 165734
rect 308394 130054 309014 165498
rect 308394 129818 308426 130054
rect 308662 129818 308746 130054
rect 308982 129818 309014 130054
rect 308394 129734 309014 129818
rect 308394 129498 308426 129734
rect 308662 129498 308746 129734
rect 308982 129498 309014 129734
rect 308394 94054 309014 129498
rect 308394 93818 308426 94054
rect 308662 93818 308746 94054
rect 308982 93818 309014 94054
rect 308394 93734 309014 93818
rect 308394 93498 308426 93734
rect 308662 93498 308746 93734
rect 308982 93498 309014 93734
rect 308394 58054 309014 93498
rect 308394 57818 308426 58054
rect 308662 57818 308746 58054
rect 308982 57818 309014 58054
rect 308394 57734 309014 57818
rect 308394 57498 308426 57734
rect 308662 57498 308746 57734
rect 308982 57498 309014 57734
rect 308394 22054 309014 57498
rect 308394 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 309014 22054
rect 308394 21734 309014 21818
rect 308394 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 309014 21734
rect 308394 -5146 309014 21498
rect 308394 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 309014 -5146
rect 308394 -5466 309014 -5382
rect 308394 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 309014 -5466
rect 308394 -7654 309014 -5702
rect 312114 710598 312734 711590
rect 312114 710362 312146 710598
rect 312382 710362 312466 710598
rect 312702 710362 312734 710598
rect 312114 710278 312734 710362
rect 312114 710042 312146 710278
rect 312382 710042 312466 710278
rect 312702 710042 312734 710278
rect 312114 673774 312734 710042
rect 312114 673538 312146 673774
rect 312382 673538 312466 673774
rect 312702 673538 312734 673774
rect 312114 673454 312734 673538
rect 312114 673218 312146 673454
rect 312382 673218 312466 673454
rect 312702 673218 312734 673454
rect 312114 637774 312734 673218
rect 312114 637538 312146 637774
rect 312382 637538 312466 637774
rect 312702 637538 312734 637774
rect 312114 637454 312734 637538
rect 312114 637218 312146 637454
rect 312382 637218 312466 637454
rect 312702 637218 312734 637454
rect 312114 601774 312734 637218
rect 312114 601538 312146 601774
rect 312382 601538 312466 601774
rect 312702 601538 312734 601774
rect 312114 601454 312734 601538
rect 312114 601218 312146 601454
rect 312382 601218 312466 601454
rect 312702 601218 312734 601454
rect 312114 565774 312734 601218
rect 312114 565538 312146 565774
rect 312382 565538 312466 565774
rect 312702 565538 312734 565774
rect 312114 565454 312734 565538
rect 312114 565218 312146 565454
rect 312382 565218 312466 565454
rect 312702 565218 312734 565454
rect 312114 529774 312734 565218
rect 312114 529538 312146 529774
rect 312382 529538 312466 529774
rect 312702 529538 312734 529774
rect 312114 529454 312734 529538
rect 312114 529218 312146 529454
rect 312382 529218 312466 529454
rect 312702 529218 312734 529454
rect 312114 493774 312734 529218
rect 312114 493538 312146 493774
rect 312382 493538 312466 493774
rect 312702 493538 312734 493774
rect 312114 493454 312734 493538
rect 312114 493218 312146 493454
rect 312382 493218 312466 493454
rect 312702 493218 312734 493454
rect 312114 457774 312734 493218
rect 312114 457538 312146 457774
rect 312382 457538 312466 457774
rect 312702 457538 312734 457774
rect 312114 457454 312734 457538
rect 312114 457218 312146 457454
rect 312382 457218 312466 457454
rect 312702 457218 312734 457454
rect 312114 421774 312734 457218
rect 312114 421538 312146 421774
rect 312382 421538 312466 421774
rect 312702 421538 312734 421774
rect 312114 421454 312734 421538
rect 312114 421218 312146 421454
rect 312382 421218 312466 421454
rect 312702 421218 312734 421454
rect 312114 385774 312734 421218
rect 312114 385538 312146 385774
rect 312382 385538 312466 385774
rect 312702 385538 312734 385774
rect 312114 385454 312734 385538
rect 312114 385218 312146 385454
rect 312382 385218 312466 385454
rect 312702 385218 312734 385454
rect 312114 349774 312734 385218
rect 312114 349538 312146 349774
rect 312382 349538 312466 349774
rect 312702 349538 312734 349774
rect 312114 349454 312734 349538
rect 312114 349218 312146 349454
rect 312382 349218 312466 349454
rect 312702 349218 312734 349454
rect 312114 313774 312734 349218
rect 312114 313538 312146 313774
rect 312382 313538 312466 313774
rect 312702 313538 312734 313774
rect 312114 313454 312734 313538
rect 312114 313218 312146 313454
rect 312382 313218 312466 313454
rect 312702 313218 312734 313454
rect 312114 277774 312734 313218
rect 312114 277538 312146 277774
rect 312382 277538 312466 277774
rect 312702 277538 312734 277774
rect 312114 277454 312734 277538
rect 312114 277218 312146 277454
rect 312382 277218 312466 277454
rect 312702 277218 312734 277454
rect 312114 241774 312734 277218
rect 312114 241538 312146 241774
rect 312382 241538 312466 241774
rect 312702 241538 312734 241774
rect 312114 241454 312734 241538
rect 312114 241218 312146 241454
rect 312382 241218 312466 241454
rect 312702 241218 312734 241454
rect 312114 205774 312734 241218
rect 312114 205538 312146 205774
rect 312382 205538 312466 205774
rect 312702 205538 312734 205774
rect 312114 205454 312734 205538
rect 312114 205218 312146 205454
rect 312382 205218 312466 205454
rect 312702 205218 312734 205454
rect 312114 169774 312734 205218
rect 312114 169538 312146 169774
rect 312382 169538 312466 169774
rect 312702 169538 312734 169774
rect 312114 169454 312734 169538
rect 312114 169218 312146 169454
rect 312382 169218 312466 169454
rect 312702 169218 312734 169454
rect 312114 133774 312734 169218
rect 312114 133538 312146 133774
rect 312382 133538 312466 133774
rect 312702 133538 312734 133774
rect 312114 133454 312734 133538
rect 312114 133218 312146 133454
rect 312382 133218 312466 133454
rect 312702 133218 312734 133454
rect 312114 97774 312734 133218
rect 312114 97538 312146 97774
rect 312382 97538 312466 97774
rect 312702 97538 312734 97774
rect 312114 97454 312734 97538
rect 312114 97218 312146 97454
rect 312382 97218 312466 97454
rect 312702 97218 312734 97454
rect 312114 61774 312734 97218
rect 312114 61538 312146 61774
rect 312382 61538 312466 61774
rect 312702 61538 312734 61774
rect 312114 61454 312734 61538
rect 312114 61218 312146 61454
rect 312382 61218 312466 61454
rect 312702 61218 312734 61454
rect 312114 25774 312734 61218
rect 312114 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 312734 25774
rect 312114 25454 312734 25538
rect 312114 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 312734 25454
rect 312114 -6106 312734 25218
rect 312114 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 312734 -6106
rect 312114 -6426 312734 -6342
rect 312114 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 312734 -6426
rect 312114 -7654 312734 -6662
rect 315834 711558 316454 711590
rect 315834 711322 315866 711558
rect 316102 711322 316186 711558
rect 316422 711322 316454 711558
rect 315834 711238 316454 711322
rect 315834 711002 315866 711238
rect 316102 711002 316186 711238
rect 316422 711002 316454 711238
rect 315834 677494 316454 711002
rect 315834 677258 315866 677494
rect 316102 677258 316186 677494
rect 316422 677258 316454 677494
rect 315834 677174 316454 677258
rect 315834 676938 315866 677174
rect 316102 676938 316186 677174
rect 316422 676938 316454 677174
rect 315834 641494 316454 676938
rect 315834 641258 315866 641494
rect 316102 641258 316186 641494
rect 316422 641258 316454 641494
rect 315834 641174 316454 641258
rect 315834 640938 315866 641174
rect 316102 640938 316186 641174
rect 316422 640938 316454 641174
rect 315834 605494 316454 640938
rect 315834 605258 315866 605494
rect 316102 605258 316186 605494
rect 316422 605258 316454 605494
rect 315834 605174 316454 605258
rect 315834 604938 315866 605174
rect 316102 604938 316186 605174
rect 316422 604938 316454 605174
rect 315834 569494 316454 604938
rect 315834 569258 315866 569494
rect 316102 569258 316186 569494
rect 316422 569258 316454 569494
rect 315834 569174 316454 569258
rect 315834 568938 315866 569174
rect 316102 568938 316186 569174
rect 316422 568938 316454 569174
rect 315834 533494 316454 568938
rect 315834 533258 315866 533494
rect 316102 533258 316186 533494
rect 316422 533258 316454 533494
rect 315834 533174 316454 533258
rect 315834 532938 315866 533174
rect 316102 532938 316186 533174
rect 316422 532938 316454 533174
rect 315834 497494 316454 532938
rect 315834 497258 315866 497494
rect 316102 497258 316186 497494
rect 316422 497258 316454 497494
rect 315834 497174 316454 497258
rect 315834 496938 315866 497174
rect 316102 496938 316186 497174
rect 316422 496938 316454 497174
rect 315834 461494 316454 496938
rect 315834 461258 315866 461494
rect 316102 461258 316186 461494
rect 316422 461258 316454 461494
rect 315834 461174 316454 461258
rect 315834 460938 315866 461174
rect 316102 460938 316186 461174
rect 316422 460938 316454 461174
rect 315834 425494 316454 460938
rect 315834 425258 315866 425494
rect 316102 425258 316186 425494
rect 316422 425258 316454 425494
rect 315834 425174 316454 425258
rect 315834 424938 315866 425174
rect 316102 424938 316186 425174
rect 316422 424938 316454 425174
rect 315834 389494 316454 424938
rect 315834 389258 315866 389494
rect 316102 389258 316186 389494
rect 316422 389258 316454 389494
rect 315834 389174 316454 389258
rect 315834 388938 315866 389174
rect 316102 388938 316186 389174
rect 316422 388938 316454 389174
rect 315834 353494 316454 388938
rect 315834 353258 315866 353494
rect 316102 353258 316186 353494
rect 316422 353258 316454 353494
rect 315834 353174 316454 353258
rect 315834 352938 315866 353174
rect 316102 352938 316186 353174
rect 316422 352938 316454 353174
rect 315834 317494 316454 352938
rect 315834 317258 315866 317494
rect 316102 317258 316186 317494
rect 316422 317258 316454 317494
rect 315834 317174 316454 317258
rect 315834 316938 315866 317174
rect 316102 316938 316186 317174
rect 316422 316938 316454 317174
rect 315834 281494 316454 316938
rect 315834 281258 315866 281494
rect 316102 281258 316186 281494
rect 316422 281258 316454 281494
rect 315834 281174 316454 281258
rect 315834 280938 315866 281174
rect 316102 280938 316186 281174
rect 316422 280938 316454 281174
rect 315834 245494 316454 280938
rect 315834 245258 315866 245494
rect 316102 245258 316186 245494
rect 316422 245258 316454 245494
rect 315834 245174 316454 245258
rect 315834 244938 315866 245174
rect 316102 244938 316186 245174
rect 316422 244938 316454 245174
rect 315834 209494 316454 244938
rect 315834 209258 315866 209494
rect 316102 209258 316186 209494
rect 316422 209258 316454 209494
rect 315834 209174 316454 209258
rect 315834 208938 315866 209174
rect 316102 208938 316186 209174
rect 316422 208938 316454 209174
rect 315834 173494 316454 208938
rect 315834 173258 315866 173494
rect 316102 173258 316186 173494
rect 316422 173258 316454 173494
rect 315834 173174 316454 173258
rect 315834 172938 315866 173174
rect 316102 172938 316186 173174
rect 316422 172938 316454 173174
rect 315834 137494 316454 172938
rect 315834 137258 315866 137494
rect 316102 137258 316186 137494
rect 316422 137258 316454 137494
rect 315834 137174 316454 137258
rect 315834 136938 315866 137174
rect 316102 136938 316186 137174
rect 316422 136938 316454 137174
rect 315834 101494 316454 136938
rect 315834 101258 315866 101494
rect 316102 101258 316186 101494
rect 316422 101258 316454 101494
rect 315834 101174 316454 101258
rect 315834 100938 315866 101174
rect 316102 100938 316186 101174
rect 316422 100938 316454 101174
rect 315834 65494 316454 100938
rect 315834 65258 315866 65494
rect 316102 65258 316186 65494
rect 316422 65258 316454 65494
rect 315834 65174 316454 65258
rect 315834 64938 315866 65174
rect 316102 64938 316186 65174
rect 316422 64938 316454 65174
rect 315834 29494 316454 64938
rect 315834 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 316454 29494
rect 315834 29174 316454 29258
rect 315834 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 316454 29174
rect 315834 -7066 316454 28938
rect 315834 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 316454 -7066
rect 315834 -7386 316454 -7302
rect 315834 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 316454 -7386
rect 315834 -7654 316454 -7622
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 329514 705798 330134 711590
rect 329514 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 330134 705798
rect 329514 705478 330134 705562
rect 329514 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 330134 705478
rect 329514 691174 330134 705242
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -1306 330134 6618
rect 329514 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 330134 -1306
rect 329514 -1626 330134 -1542
rect 329514 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 330134 -1626
rect 329514 -7654 330134 -1862
rect 333234 706758 333854 711590
rect 333234 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 333854 706758
rect 333234 706438 333854 706522
rect 333234 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 333854 706438
rect 333234 694894 333854 706202
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -2266 333854 10338
rect 333234 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 333854 -2266
rect 333234 -2586 333854 -2502
rect 333234 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 333854 -2586
rect 333234 -7654 333854 -2822
rect 336954 707718 337574 711590
rect 336954 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 337574 707718
rect 336954 707398 337574 707482
rect 336954 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 337574 707398
rect 336954 698614 337574 707162
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 336954 -3226 337574 14058
rect 336954 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 337574 -3226
rect 336954 -3546 337574 -3462
rect 336954 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 337574 -3546
rect 336954 -7654 337574 -3782
rect 340674 708678 341294 711590
rect 340674 708442 340706 708678
rect 340942 708442 341026 708678
rect 341262 708442 341294 708678
rect 340674 708358 341294 708442
rect 340674 708122 340706 708358
rect 340942 708122 341026 708358
rect 341262 708122 341294 708358
rect 340674 666334 341294 708122
rect 340674 666098 340706 666334
rect 340942 666098 341026 666334
rect 341262 666098 341294 666334
rect 340674 666014 341294 666098
rect 340674 665778 340706 666014
rect 340942 665778 341026 666014
rect 341262 665778 341294 666014
rect 340674 630334 341294 665778
rect 340674 630098 340706 630334
rect 340942 630098 341026 630334
rect 341262 630098 341294 630334
rect 340674 630014 341294 630098
rect 340674 629778 340706 630014
rect 340942 629778 341026 630014
rect 341262 629778 341294 630014
rect 340674 594334 341294 629778
rect 340674 594098 340706 594334
rect 340942 594098 341026 594334
rect 341262 594098 341294 594334
rect 340674 594014 341294 594098
rect 340674 593778 340706 594014
rect 340942 593778 341026 594014
rect 341262 593778 341294 594014
rect 340674 558334 341294 593778
rect 340674 558098 340706 558334
rect 340942 558098 341026 558334
rect 341262 558098 341294 558334
rect 340674 558014 341294 558098
rect 340674 557778 340706 558014
rect 340942 557778 341026 558014
rect 341262 557778 341294 558014
rect 340674 522334 341294 557778
rect 340674 522098 340706 522334
rect 340942 522098 341026 522334
rect 341262 522098 341294 522334
rect 340674 522014 341294 522098
rect 340674 521778 340706 522014
rect 340942 521778 341026 522014
rect 341262 521778 341294 522014
rect 340674 486334 341294 521778
rect 340674 486098 340706 486334
rect 340942 486098 341026 486334
rect 341262 486098 341294 486334
rect 340674 486014 341294 486098
rect 340674 485778 340706 486014
rect 340942 485778 341026 486014
rect 341262 485778 341294 486014
rect 340674 450334 341294 485778
rect 340674 450098 340706 450334
rect 340942 450098 341026 450334
rect 341262 450098 341294 450334
rect 340674 450014 341294 450098
rect 340674 449778 340706 450014
rect 340942 449778 341026 450014
rect 341262 449778 341294 450014
rect 340674 414334 341294 449778
rect 340674 414098 340706 414334
rect 340942 414098 341026 414334
rect 341262 414098 341294 414334
rect 340674 414014 341294 414098
rect 340674 413778 340706 414014
rect 340942 413778 341026 414014
rect 341262 413778 341294 414014
rect 340674 378334 341294 413778
rect 340674 378098 340706 378334
rect 340942 378098 341026 378334
rect 341262 378098 341294 378334
rect 340674 378014 341294 378098
rect 340674 377778 340706 378014
rect 340942 377778 341026 378014
rect 341262 377778 341294 378014
rect 340674 342334 341294 377778
rect 340674 342098 340706 342334
rect 340942 342098 341026 342334
rect 341262 342098 341294 342334
rect 340674 342014 341294 342098
rect 340674 341778 340706 342014
rect 340942 341778 341026 342014
rect 341262 341778 341294 342014
rect 340674 306334 341294 341778
rect 340674 306098 340706 306334
rect 340942 306098 341026 306334
rect 341262 306098 341294 306334
rect 340674 306014 341294 306098
rect 340674 305778 340706 306014
rect 340942 305778 341026 306014
rect 341262 305778 341294 306014
rect 340674 270334 341294 305778
rect 340674 270098 340706 270334
rect 340942 270098 341026 270334
rect 341262 270098 341294 270334
rect 340674 270014 341294 270098
rect 340674 269778 340706 270014
rect 340942 269778 341026 270014
rect 341262 269778 341294 270014
rect 340674 234334 341294 269778
rect 340674 234098 340706 234334
rect 340942 234098 341026 234334
rect 341262 234098 341294 234334
rect 340674 234014 341294 234098
rect 340674 233778 340706 234014
rect 340942 233778 341026 234014
rect 341262 233778 341294 234014
rect 340674 198334 341294 233778
rect 340674 198098 340706 198334
rect 340942 198098 341026 198334
rect 341262 198098 341294 198334
rect 340674 198014 341294 198098
rect 340674 197778 340706 198014
rect 340942 197778 341026 198014
rect 341262 197778 341294 198014
rect 340674 162334 341294 197778
rect 340674 162098 340706 162334
rect 340942 162098 341026 162334
rect 341262 162098 341294 162334
rect 340674 162014 341294 162098
rect 340674 161778 340706 162014
rect 340942 161778 341026 162014
rect 341262 161778 341294 162014
rect 340674 126334 341294 161778
rect 340674 126098 340706 126334
rect 340942 126098 341026 126334
rect 341262 126098 341294 126334
rect 340674 126014 341294 126098
rect 340674 125778 340706 126014
rect 340942 125778 341026 126014
rect 341262 125778 341294 126014
rect 340674 90334 341294 125778
rect 340674 90098 340706 90334
rect 340942 90098 341026 90334
rect 341262 90098 341294 90334
rect 340674 90014 341294 90098
rect 340674 89778 340706 90014
rect 340942 89778 341026 90014
rect 341262 89778 341294 90014
rect 340674 54334 341294 89778
rect 340674 54098 340706 54334
rect 340942 54098 341026 54334
rect 341262 54098 341294 54334
rect 340674 54014 341294 54098
rect 340674 53778 340706 54014
rect 340942 53778 341026 54014
rect 341262 53778 341294 54014
rect 340674 18334 341294 53778
rect 340674 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 341294 18334
rect 340674 18014 341294 18098
rect 340674 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 341294 18014
rect 340674 -4186 341294 17778
rect 340674 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 341294 -4186
rect 340674 -4506 341294 -4422
rect 340674 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 341294 -4506
rect 340674 -7654 341294 -4742
rect 344394 709638 345014 711590
rect 344394 709402 344426 709638
rect 344662 709402 344746 709638
rect 344982 709402 345014 709638
rect 344394 709318 345014 709402
rect 344394 709082 344426 709318
rect 344662 709082 344746 709318
rect 344982 709082 345014 709318
rect 344394 670054 345014 709082
rect 344394 669818 344426 670054
rect 344662 669818 344746 670054
rect 344982 669818 345014 670054
rect 344394 669734 345014 669818
rect 344394 669498 344426 669734
rect 344662 669498 344746 669734
rect 344982 669498 345014 669734
rect 344394 634054 345014 669498
rect 344394 633818 344426 634054
rect 344662 633818 344746 634054
rect 344982 633818 345014 634054
rect 344394 633734 345014 633818
rect 344394 633498 344426 633734
rect 344662 633498 344746 633734
rect 344982 633498 345014 633734
rect 344394 598054 345014 633498
rect 344394 597818 344426 598054
rect 344662 597818 344746 598054
rect 344982 597818 345014 598054
rect 344394 597734 345014 597818
rect 344394 597498 344426 597734
rect 344662 597498 344746 597734
rect 344982 597498 345014 597734
rect 344394 562054 345014 597498
rect 344394 561818 344426 562054
rect 344662 561818 344746 562054
rect 344982 561818 345014 562054
rect 344394 561734 345014 561818
rect 344394 561498 344426 561734
rect 344662 561498 344746 561734
rect 344982 561498 345014 561734
rect 344394 526054 345014 561498
rect 344394 525818 344426 526054
rect 344662 525818 344746 526054
rect 344982 525818 345014 526054
rect 344394 525734 345014 525818
rect 344394 525498 344426 525734
rect 344662 525498 344746 525734
rect 344982 525498 345014 525734
rect 344394 490054 345014 525498
rect 344394 489818 344426 490054
rect 344662 489818 344746 490054
rect 344982 489818 345014 490054
rect 344394 489734 345014 489818
rect 344394 489498 344426 489734
rect 344662 489498 344746 489734
rect 344982 489498 345014 489734
rect 344394 454054 345014 489498
rect 344394 453818 344426 454054
rect 344662 453818 344746 454054
rect 344982 453818 345014 454054
rect 344394 453734 345014 453818
rect 344394 453498 344426 453734
rect 344662 453498 344746 453734
rect 344982 453498 345014 453734
rect 344394 418054 345014 453498
rect 344394 417818 344426 418054
rect 344662 417818 344746 418054
rect 344982 417818 345014 418054
rect 344394 417734 345014 417818
rect 344394 417498 344426 417734
rect 344662 417498 344746 417734
rect 344982 417498 345014 417734
rect 344394 382054 345014 417498
rect 344394 381818 344426 382054
rect 344662 381818 344746 382054
rect 344982 381818 345014 382054
rect 344394 381734 345014 381818
rect 344394 381498 344426 381734
rect 344662 381498 344746 381734
rect 344982 381498 345014 381734
rect 344394 346054 345014 381498
rect 344394 345818 344426 346054
rect 344662 345818 344746 346054
rect 344982 345818 345014 346054
rect 344394 345734 345014 345818
rect 344394 345498 344426 345734
rect 344662 345498 344746 345734
rect 344982 345498 345014 345734
rect 344394 310054 345014 345498
rect 344394 309818 344426 310054
rect 344662 309818 344746 310054
rect 344982 309818 345014 310054
rect 344394 309734 345014 309818
rect 344394 309498 344426 309734
rect 344662 309498 344746 309734
rect 344982 309498 345014 309734
rect 344394 274054 345014 309498
rect 344394 273818 344426 274054
rect 344662 273818 344746 274054
rect 344982 273818 345014 274054
rect 344394 273734 345014 273818
rect 344394 273498 344426 273734
rect 344662 273498 344746 273734
rect 344982 273498 345014 273734
rect 344394 238054 345014 273498
rect 344394 237818 344426 238054
rect 344662 237818 344746 238054
rect 344982 237818 345014 238054
rect 344394 237734 345014 237818
rect 344394 237498 344426 237734
rect 344662 237498 344746 237734
rect 344982 237498 345014 237734
rect 344394 202054 345014 237498
rect 344394 201818 344426 202054
rect 344662 201818 344746 202054
rect 344982 201818 345014 202054
rect 344394 201734 345014 201818
rect 344394 201498 344426 201734
rect 344662 201498 344746 201734
rect 344982 201498 345014 201734
rect 344394 166054 345014 201498
rect 344394 165818 344426 166054
rect 344662 165818 344746 166054
rect 344982 165818 345014 166054
rect 344394 165734 345014 165818
rect 344394 165498 344426 165734
rect 344662 165498 344746 165734
rect 344982 165498 345014 165734
rect 344394 130054 345014 165498
rect 344394 129818 344426 130054
rect 344662 129818 344746 130054
rect 344982 129818 345014 130054
rect 344394 129734 345014 129818
rect 344394 129498 344426 129734
rect 344662 129498 344746 129734
rect 344982 129498 345014 129734
rect 344394 94054 345014 129498
rect 344394 93818 344426 94054
rect 344662 93818 344746 94054
rect 344982 93818 345014 94054
rect 344394 93734 345014 93818
rect 344394 93498 344426 93734
rect 344662 93498 344746 93734
rect 344982 93498 345014 93734
rect 344394 58054 345014 93498
rect 344394 57818 344426 58054
rect 344662 57818 344746 58054
rect 344982 57818 345014 58054
rect 344394 57734 345014 57818
rect 344394 57498 344426 57734
rect 344662 57498 344746 57734
rect 344982 57498 345014 57734
rect 344394 22054 345014 57498
rect 344394 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 345014 22054
rect 344394 21734 345014 21818
rect 344394 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 345014 21734
rect 344394 -5146 345014 21498
rect 344394 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 345014 -5146
rect 344394 -5466 345014 -5382
rect 344394 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 345014 -5466
rect 344394 -7654 345014 -5702
rect 348114 710598 348734 711590
rect 348114 710362 348146 710598
rect 348382 710362 348466 710598
rect 348702 710362 348734 710598
rect 348114 710278 348734 710362
rect 348114 710042 348146 710278
rect 348382 710042 348466 710278
rect 348702 710042 348734 710278
rect 348114 673774 348734 710042
rect 348114 673538 348146 673774
rect 348382 673538 348466 673774
rect 348702 673538 348734 673774
rect 348114 673454 348734 673538
rect 348114 673218 348146 673454
rect 348382 673218 348466 673454
rect 348702 673218 348734 673454
rect 348114 637774 348734 673218
rect 348114 637538 348146 637774
rect 348382 637538 348466 637774
rect 348702 637538 348734 637774
rect 348114 637454 348734 637538
rect 348114 637218 348146 637454
rect 348382 637218 348466 637454
rect 348702 637218 348734 637454
rect 348114 601774 348734 637218
rect 348114 601538 348146 601774
rect 348382 601538 348466 601774
rect 348702 601538 348734 601774
rect 348114 601454 348734 601538
rect 348114 601218 348146 601454
rect 348382 601218 348466 601454
rect 348702 601218 348734 601454
rect 348114 565774 348734 601218
rect 348114 565538 348146 565774
rect 348382 565538 348466 565774
rect 348702 565538 348734 565774
rect 348114 565454 348734 565538
rect 348114 565218 348146 565454
rect 348382 565218 348466 565454
rect 348702 565218 348734 565454
rect 348114 529774 348734 565218
rect 348114 529538 348146 529774
rect 348382 529538 348466 529774
rect 348702 529538 348734 529774
rect 348114 529454 348734 529538
rect 348114 529218 348146 529454
rect 348382 529218 348466 529454
rect 348702 529218 348734 529454
rect 348114 493774 348734 529218
rect 348114 493538 348146 493774
rect 348382 493538 348466 493774
rect 348702 493538 348734 493774
rect 348114 493454 348734 493538
rect 348114 493218 348146 493454
rect 348382 493218 348466 493454
rect 348702 493218 348734 493454
rect 348114 457774 348734 493218
rect 348114 457538 348146 457774
rect 348382 457538 348466 457774
rect 348702 457538 348734 457774
rect 348114 457454 348734 457538
rect 348114 457218 348146 457454
rect 348382 457218 348466 457454
rect 348702 457218 348734 457454
rect 348114 421774 348734 457218
rect 348114 421538 348146 421774
rect 348382 421538 348466 421774
rect 348702 421538 348734 421774
rect 348114 421454 348734 421538
rect 348114 421218 348146 421454
rect 348382 421218 348466 421454
rect 348702 421218 348734 421454
rect 348114 385774 348734 421218
rect 348114 385538 348146 385774
rect 348382 385538 348466 385774
rect 348702 385538 348734 385774
rect 348114 385454 348734 385538
rect 348114 385218 348146 385454
rect 348382 385218 348466 385454
rect 348702 385218 348734 385454
rect 348114 349774 348734 385218
rect 348114 349538 348146 349774
rect 348382 349538 348466 349774
rect 348702 349538 348734 349774
rect 348114 349454 348734 349538
rect 348114 349218 348146 349454
rect 348382 349218 348466 349454
rect 348702 349218 348734 349454
rect 348114 313774 348734 349218
rect 348114 313538 348146 313774
rect 348382 313538 348466 313774
rect 348702 313538 348734 313774
rect 348114 313454 348734 313538
rect 348114 313218 348146 313454
rect 348382 313218 348466 313454
rect 348702 313218 348734 313454
rect 348114 277774 348734 313218
rect 348114 277538 348146 277774
rect 348382 277538 348466 277774
rect 348702 277538 348734 277774
rect 348114 277454 348734 277538
rect 348114 277218 348146 277454
rect 348382 277218 348466 277454
rect 348702 277218 348734 277454
rect 348114 241774 348734 277218
rect 348114 241538 348146 241774
rect 348382 241538 348466 241774
rect 348702 241538 348734 241774
rect 348114 241454 348734 241538
rect 348114 241218 348146 241454
rect 348382 241218 348466 241454
rect 348702 241218 348734 241454
rect 348114 205774 348734 241218
rect 348114 205538 348146 205774
rect 348382 205538 348466 205774
rect 348702 205538 348734 205774
rect 348114 205454 348734 205538
rect 348114 205218 348146 205454
rect 348382 205218 348466 205454
rect 348702 205218 348734 205454
rect 348114 169774 348734 205218
rect 348114 169538 348146 169774
rect 348382 169538 348466 169774
rect 348702 169538 348734 169774
rect 348114 169454 348734 169538
rect 348114 169218 348146 169454
rect 348382 169218 348466 169454
rect 348702 169218 348734 169454
rect 348114 133774 348734 169218
rect 348114 133538 348146 133774
rect 348382 133538 348466 133774
rect 348702 133538 348734 133774
rect 348114 133454 348734 133538
rect 348114 133218 348146 133454
rect 348382 133218 348466 133454
rect 348702 133218 348734 133454
rect 348114 97774 348734 133218
rect 348114 97538 348146 97774
rect 348382 97538 348466 97774
rect 348702 97538 348734 97774
rect 348114 97454 348734 97538
rect 348114 97218 348146 97454
rect 348382 97218 348466 97454
rect 348702 97218 348734 97454
rect 348114 61774 348734 97218
rect 348114 61538 348146 61774
rect 348382 61538 348466 61774
rect 348702 61538 348734 61774
rect 348114 61454 348734 61538
rect 348114 61218 348146 61454
rect 348382 61218 348466 61454
rect 348702 61218 348734 61454
rect 348114 25774 348734 61218
rect 348114 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 348734 25774
rect 348114 25454 348734 25538
rect 348114 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 348734 25454
rect 348114 -6106 348734 25218
rect 348114 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 348734 -6106
rect 348114 -6426 348734 -6342
rect 348114 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 348734 -6426
rect 348114 -7654 348734 -6662
rect 351834 711558 352454 711590
rect 351834 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 352454 711558
rect 351834 711238 352454 711322
rect 351834 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 352454 711238
rect 351834 677494 352454 711002
rect 351834 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 352454 677494
rect 351834 677174 352454 677258
rect 351834 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 352454 677174
rect 351834 641494 352454 676938
rect 351834 641258 351866 641494
rect 352102 641258 352186 641494
rect 352422 641258 352454 641494
rect 351834 641174 352454 641258
rect 351834 640938 351866 641174
rect 352102 640938 352186 641174
rect 352422 640938 352454 641174
rect 351834 605494 352454 640938
rect 351834 605258 351866 605494
rect 352102 605258 352186 605494
rect 352422 605258 352454 605494
rect 351834 605174 352454 605258
rect 351834 604938 351866 605174
rect 352102 604938 352186 605174
rect 352422 604938 352454 605174
rect 351834 569494 352454 604938
rect 351834 569258 351866 569494
rect 352102 569258 352186 569494
rect 352422 569258 352454 569494
rect 351834 569174 352454 569258
rect 351834 568938 351866 569174
rect 352102 568938 352186 569174
rect 352422 568938 352454 569174
rect 351834 533494 352454 568938
rect 351834 533258 351866 533494
rect 352102 533258 352186 533494
rect 352422 533258 352454 533494
rect 351834 533174 352454 533258
rect 351834 532938 351866 533174
rect 352102 532938 352186 533174
rect 352422 532938 352454 533174
rect 351834 497494 352454 532938
rect 351834 497258 351866 497494
rect 352102 497258 352186 497494
rect 352422 497258 352454 497494
rect 351834 497174 352454 497258
rect 351834 496938 351866 497174
rect 352102 496938 352186 497174
rect 352422 496938 352454 497174
rect 351834 461494 352454 496938
rect 351834 461258 351866 461494
rect 352102 461258 352186 461494
rect 352422 461258 352454 461494
rect 351834 461174 352454 461258
rect 351834 460938 351866 461174
rect 352102 460938 352186 461174
rect 352422 460938 352454 461174
rect 351834 425494 352454 460938
rect 351834 425258 351866 425494
rect 352102 425258 352186 425494
rect 352422 425258 352454 425494
rect 351834 425174 352454 425258
rect 351834 424938 351866 425174
rect 352102 424938 352186 425174
rect 352422 424938 352454 425174
rect 351834 389494 352454 424938
rect 351834 389258 351866 389494
rect 352102 389258 352186 389494
rect 352422 389258 352454 389494
rect 351834 389174 352454 389258
rect 351834 388938 351866 389174
rect 352102 388938 352186 389174
rect 352422 388938 352454 389174
rect 351834 353494 352454 388938
rect 351834 353258 351866 353494
rect 352102 353258 352186 353494
rect 352422 353258 352454 353494
rect 351834 353174 352454 353258
rect 351834 352938 351866 353174
rect 352102 352938 352186 353174
rect 352422 352938 352454 353174
rect 351834 317494 352454 352938
rect 351834 317258 351866 317494
rect 352102 317258 352186 317494
rect 352422 317258 352454 317494
rect 351834 317174 352454 317258
rect 351834 316938 351866 317174
rect 352102 316938 352186 317174
rect 352422 316938 352454 317174
rect 351834 281494 352454 316938
rect 351834 281258 351866 281494
rect 352102 281258 352186 281494
rect 352422 281258 352454 281494
rect 351834 281174 352454 281258
rect 351834 280938 351866 281174
rect 352102 280938 352186 281174
rect 352422 280938 352454 281174
rect 351834 245494 352454 280938
rect 351834 245258 351866 245494
rect 352102 245258 352186 245494
rect 352422 245258 352454 245494
rect 351834 245174 352454 245258
rect 351834 244938 351866 245174
rect 352102 244938 352186 245174
rect 352422 244938 352454 245174
rect 351834 209494 352454 244938
rect 351834 209258 351866 209494
rect 352102 209258 352186 209494
rect 352422 209258 352454 209494
rect 351834 209174 352454 209258
rect 351834 208938 351866 209174
rect 352102 208938 352186 209174
rect 352422 208938 352454 209174
rect 351834 173494 352454 208938
rect 351834 173258 351866 173494
rect 352102 173258 352186 173494
rect 352422 173258 352454 173494
rect 351834 173174 352454 173258
rect 351834 172938 351866 173174
rect 352102 172938 352186 173174
rect 352422 172938 352454 173174
rect 351834 137494 352454 172938
rect 351834 137258 351866 137494
rect 352102 137258 352186 137494
rect 352422 137258 352454 137494
rect 351834 137174 352454 137258
rect 351834 136938 351866 137174
rect 352102 136938 352186 137174
rect 352422 136938 352454 137174
rect 351834 101494 352454 136938
rect 351834 101258 351866 101494
rect 352102 101258 352186 101494
rect 352422 101258 352454 101494
rect 351834 101174 352454 101258
rect 351834 100938 351866 101174
rect 352102 100938 352186 101174
rect 352422 100938 352454 101174
rect 351834 65494 352454 100938
rect 351834 65258 351866 65494
rect 352102 65258 352186 65494
rect 352422 65258 352454 65494
rect 351834 65174 352454 65258
rect 351834 64938 351866 65174
rect 352102 64938 352186 65174
rect 352422 64938 352454 65174
rect 351834 29494 352454 64938
rect 351834 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 352454 29494
rect 351834 29174 352454 29258
rect 351834 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 352454 29174
rect 351834 -7066 352454 28938
rect 351834 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 352454 -7066
rect 351834 -7386 352454 -7302
rect 351834 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 352454 -7386
rect 351834 -7654 352454 -7622
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 365514 705798 366134 711590
rect 365514 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 366134 705798
rect 365514 705478 366134 705562
rect 365514 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 366134 705478
rect 365514 691174 366134 705242
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -1306 366134 6618
rect 365514 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 366134 -1306
rect 365514 -1626 366134 -1542
rect 365514 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 366134 -1626
rect 365514 -7654 366134 -1862
rect 369234 706758 369854 711590
rect 369234 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 369854 706758
rect 369234 706438 369854 706522
rect 369234 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 369854 706438
rect 369234 694894 369854 706202
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -2266 369854 10338
rect 369234 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 369854 -2266
rect 369234 -2586 369854 -2502
rect 369234 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 369854 -2586
rect 369234 -7654 369854 -2822
rect 372954 707718 373574 711590
rect 372954 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 373574 707718
rect 372954 707398 373574 707482
rect 372954 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 373574 707398
rect 372954 698614 373574 707162
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 372954 -3226 373574 14058
rect 372954 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 373574 -3226
rect 372954 -3546 373574 -3462
rect 372954 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 373574 -3546
rect 372954 -7654 373574 -3782
rect 376674 708678 377294 711590
rect 376674 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 377294 708678
rect 376674 708358 377294 708442
rect 376674 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 377294 708358
rect 376674 666334 377294 708122
rect 376674 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 377294 666334
rect 376674 666014 377294 666098
rect 376674 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 377294 666014
rect 376674 630334 377294 665778
rect 376674 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 377294 630334
rect 376674 630014 377294 630098
rect 376674 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 377294 630014
rect 376674 594334 377294 629778
rect 376674 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 377294 594334
rect 376674 594014 377294 594098
rect 376674 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 377294 594014
rect 376674 558334 377294 593778
rect 376674 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 377294 558334
rect 376674 558014 377294 558098
rect 376674 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 377294 558014
rect 376674 522334 377294 557778
rect 376674 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 377294 522334
rect 376674 522014 377294 522098
rect 376674 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 377294 522014
rect 376674 486334 377294 521778
rect 376674 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 377294 486334
rect 376674 486014 377294 486098
rect 376674 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 377294 486014
rect 376674 450334 377294 485778
rect 376674 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 377294 450334
rect 376674 450014 377294 450098
rect 376674 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 377294 450014
rect 376674 414334 377294 449778
rect 376674 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 377294 414334
rect 376674 414014 377294 414098
rect 376674 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 377294 414014
rect 376674 378334 377294 413778
rect 376674 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 377294 378334
rect 376674 378014 377294 378098
rect 376674 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 377294 378014
rect 376674 342334 377294 377778
rect 376674 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 377294 342334
rect 376674 342014 377294 342098
rect 376674 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 377294 342014
rect 376674 306334 377294 341778
rect 376674 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 377294 306334
rect 376674 306014 377294 306098
rect 376674 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 377294 306014
rect 376674 270334 377294 305778
rect 376674 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 377294 270334
rect 376674 270014 377294 270098
rect 376674 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 377294 270014
rect 376674 234334 377294 269778
rect 376674 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 377294 234334
rect 376674 234014 377294 234098
rect 376674 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 377294 234014
rect 376674 198334 377294 233778
rect 376674 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 377294 198334
rect 376674 198014 377294 198098
rect 376674 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 377294 198014
rect 376674 162334 377294 197778
rect 376674 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 377294 162334
rect 376674 162014 377294 162098
rect 376674 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 377294 162014
rect 376674 126334 377294 161778
rect 376674 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 377294 126334
rect 376674 126014 377294 126098
rect 376674 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 377294 126014
rect 376674 90334 377294 125778
rect 376674 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 377294 90334
rect 376674 90014 377294 90098
rect 376674 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 377294 90014
rect 376674 54334 377294 89778
rect 376674 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 377294 54334
rect 376674 54014 377294 54098
rect 376674 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 377294 54014
rect 376674 18334 377294 53778
rect 376674 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 377294 18334
rect 376674 18014 377294 18098
rect 376674 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 377294 18014
rect 376674 -4186 377294 17778
rect 376674 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 377294 -4186
rect 376674 -4506 377294 -4422
rect 376674 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 377294 -4506
rect 376674 -7654 377294 -4742
rect 380394 709638 381014 711590
rect 380394 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 381014 709638
rect 380394 709318 381014 709402
rect 380394 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 381014 709318
rect 380394 670054 381014 709082
rect 380394 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 381014 670054
rect 380394 669734 381014 669818
rect 380394 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 381014 669734
rect 380394 634054 381014 669498
rect 380394 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 381014 634054
rect 380394 633734 381014 633818
rect 380394 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 381014 633734
rect 380394 598054 381014 633498
rect 380394 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 381014 598054
rect 380394 597734 381014 597818
rect 380394 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 381014 597734
rect 380394 562054 381014 597498
rect 380394 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 381014 562054
rect 380394 561734 381014 561818
rect 380394 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 381014 561734
rect 380394 526054 381014 561498
rect 380394 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 381014 526054
rect 380394 525734 381014 525818
rect 380394 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 381014 525734
rect 380394 490054 381014 525498
rect 380394 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 381014 490054
rect 380394 489734 381014 489818
rect 380394 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 381014 489734
rect 380394 454054 381014 489498
rect 380394 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 381014 454054
rect 380394 453734 381014 453818
rect 380394 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 381014 453734
rect 380394 418054 381014 453498
rect 380394 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 381014 418054
rect 380394 417734 381014 417818
rect 380394 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 381014 417734
rect 380394 382054 381014 417498
rect 380394 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 381014 382054
rect 380394 381734 381014 381818
rect 380394 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 381014 381734
rect 380394 346054 381014 381498
rect 380394 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 381014 346054
rect 380394 345734 381014 345818
rect 380394 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 381014 345734
rect 380394 310054 381014 345498
rect 380394 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 381014 310054
rect 380394 309734 381014 309818
rect 380394 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 381014 309734
rect 380394 274054 381014 309498
rect 380394 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 381014 274054
rect 380394 273734 381014 273818
rect 380394 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 381014 273734
rect 380394 238054 381014 273498
rect 380394 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 381014 238054
rect 380394 237734 381014 237818
rect 380394 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 381014 237734
rect 380394 202054 381014 237498
rect 380394 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 381014 202054
rect 380394 201734 381014 201818
rect 380394 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 381014 201734
rect 380394 166054 381014 201498
rect 380394 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 381014 166054
rect 380394 165734 381014 165818
rect 380394 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 381014 165734
rect 380394 130054 381014 165498
rect 380394 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 381014 130054
rect 380394 129734 381014 129818
rect 380394 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 381014 129734
rect 380394 94054 381014 129498
rect 380394 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 381014 94054
rect 380394 93734 381014 93818
rect 380394 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 381014 93734
rect 380394 58054 381014 93498
rect 380394 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 381014 58054
rect 380394 57734 381014 57818
rect 380394 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 381014 57734
rect 380394 22054 381014 57498
rect 380394 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 381014 22054
rect 380394 21734 381014 21818
rect 380394 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 381014 21734
rect 380394 -5146 381014 21498
rect 380394 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 381014 -5146
rect 380394 -5466 381014 -5382
rect 380394 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 381014 -5466
rect 380394 -7654 381014 -5702
rect 384114 710598 384734 711590
rect 384114 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 384734 710598
rect 384114 710278 384734 710362
rect 384114 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 384734 710278
rect 384114 673774 384734 710042
rect 384114 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 384734 673774
rect 384114 673454 384734 673538
rect 384114 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 384734 673454
rect 384114 637774 384734 673218
rect 384114 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 384734 637774
rect 384114 637454 384734 637538
rect 384114 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 384734 637454
rect 384114 601774 384734 637218
rect 384114 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 384734 601774
rect 384114 601454 384734 601538
rect 384114 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 384734 601454
rect 384114 565774 384734 601218
rect 384114 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 384734 565774
rect 384114 565454 384734 565538
rect 384114 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 384734 565454
rect 384114 529774 384734 565218
rect 384114 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 384734 529774
rect 384114 529454 384734 529538
rect 384114 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 384734 529454
rect 384114 493774 384734 529218
rect 384114 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 384734 493774
rect 384114 493454 384734 493538
rect 384114 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 384734 493454
rect 384114 457774 384734 493218
rect 384114 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 384734 457774
rect 384114 457454 384734 457538
rect 384114 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 384734 457454
rect 384114 421774 384734 457218
rect 384114 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 384734 421774
rect 384114 421454 384734 421538
rect 384114 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 384734 421454
rect 384114 385774 384734 421218
rect 384114 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 384734 385774
rect 384114 385454 384734 385538
rect 384114 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 384734 385454
rect 384114 349774 384734 385218
rect 384114 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 384734 349774
rect 384114 349454 384734 349538
rect 384114 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 384734 349454
rect 384114 313774 384734 349218
rect 384114 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 384734 313774
rect 384114 313454 384734 313538
rect 384114 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 384734 313454
rect 384114 277774 384734 313218
rect 384114 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 384734 277774
rect 384114 277454 384734 277538
rect 384114 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 384734 277454
rect 384114 241774 384734 277218
rect 384114 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 384734 241774
rect 384114 241454 384734 241538
rect 384114 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 384734 241454
rect 384114 205774 384734 241218
rect 384114 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 384734 205774
rect 384114 205454 384734 205538
rect 384114 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 384734 205454
rect 384114 169774 384734 205218
rect 384114 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 384734 169774
rect 384114 169454 384734 169538
rect 384114 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 384734 169454
rect 384114 133774 384734 169218
rect 384114 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 384734 133774
rect 384114 133454 384734 133538
rect 384114 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 384734 133454
rect 384114 97774 384734 133218
rect 384114 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 384734 97774
rect 384114 97454 384734 97538
rect 384114 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 384734 97454
rect 384114 61774 384734 97218
rect 384114 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 384734 61774
rect 384114 61454 384734 61538
rect 384114 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 384734 61454
rect 384114 25774 384734 61218
rect 384114 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 384734 25774
rect 384114 25454 384734 25538
rect 384114 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 384734 25454
rect 384114 -6106 384734 25218
rect 384114 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 384734 -6106
rect 384114 -6426 384734 -6342
rect 384114 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 384734 -6426
rect 384114 -7654 384734 -6662
rect 387834 711558 388454 711590
rect 387834 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 388454 711558
rect 387834 711238 388454 711322
rect 387834 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 388454 711238
rect 387834 677494 388454 711002
rect 387834 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 388454 677494
rect 387834 677174 388454 677258
rect 387834 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 388454 677174
rect 387834 641494 388454 676938
rect 387834 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 388454 641494
rect 387834 641174 388454 641258
rect 387834 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 388454 641174
rect 387834 605494 388454 640938
rect 387834 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 388454 605494
rect 387834 605174 388454 605258
rect 387834 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 388454 605174
rect 387834 569494 388454 604938
rect 387834 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 388454 569494
rect 387834 569174 388454 569258
rect 387834 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 388454 569174
rect 387834 533494 388454 568938
rect 387834 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 388454 533494
rect 387834 533174 388454 533258
rect 387834 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 388454 533174
rect 387834 497494 388454 532938
rect 387834 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 388454 497494
rect 387834 497174 388454 497258
rect 387834 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 388454 497174
rect 387834 461494 388454 496938
rect 387834 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 388454 461494
rect 387834 461174 388454 461258
rect 387834 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 388454 461174
rect 387834 425494 388454 460938
rect 387834 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 388454 425494
rect 387834 425174 388454 425258
rect 387834 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 388454 425174
rect 387834 389494 388454 424938
rect 387834 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 388454 389494
rect 387834 389174 388454 389258
rect 387834 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 388454 389174
rect 387834 353494 388454 388938
rect 387834 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 388454 353494
rect 387834 353174 388454 353258
rect 387834 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 388454 353174
rect 387834 317494 388454 352938
rect 387834 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 388454 317494
rect 387834 317174 388454 317258
rect 387834 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 388454 317174
rect 387834 281494 388454 316938
rect 387834 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 388454 281494
rect 387834 281174 388454 281258
rect 387834 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 388454 281174
rect 387834 245494 388454 280938
rect 387834 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 388454 245494
rect 387834 245174 388454 245258
rect 387834 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 388454 245174
rect 387834 209494 388454 244938
rect 387834 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 388454 209494
rect 387834 209174 388454 209258
rect 387834 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 388454 209174
rect 387834 173494 388454 208938
rect 387834 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 388454 173494
rect 387834 173174 388454 173258
rect 387834 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 388454 173174
rect 387834 137494 388454 172938
rect 387834 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 388454 137494
rect 387834 137174 388454 137258
rect 387834 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 388454 137174
rect 387834 101494 388454 136938
rect 387834 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 388454 101494
rect 387834 101174 388454 101258
rect 387834 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 388454 101174
rect 387834 65494 388454 100938
rect 387834 65258 387866 65494
rect 388102 65258 388186 65494
rect 388422 65258 388454 65494
rect 387834 65174 388454 65258
rect 387834 64938 387866 65174
rect 388102 64938 388186 65174
rect 388422 64938 388454 65174
rect 387834 29494 388454 64938
rect 387834 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 388454 29494
rect 387834 29174 388454 29258
rect 387834 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 388454 29174
rect 387834 -7066 388454 28938
rect 387834 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 388454 -7066
rect 387834 -7386 388454 -7302
rect 387834 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 388454 -7386
rect 387834 -7654 388454 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 401514 705798 402134 711590
rect 401514 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 402134 705798
rect 401514 705478 402134 705562
rect 401514 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 402134 705478
rect 401514 691174 402134 705242
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -1306 402134 6618
rect 401514 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 402134 -1306
rect 401514 -1626 402134 -1542
rect 401514 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 402134 -1626
rect 401514 -7654 402134 -1862
rect 405234 706758 405854 711590
rect 405234 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 405854 706758
rect 405234 706438 405854 706522
rect 405234 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 405854 706438
rect 405234 694894 405854 706202
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -2266 405854 10338
rect 405234 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 405854 -2266
rect 405234 -2586 405854 -2502
rect 405234 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 405854 -2586
rect 405234 -7654 405854 -2822
rect 408954 707718 409574 711590
rect 408954 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 409574 707718
rect 408954 707398 409574 707482
rect 408954 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 409574 707398
rect 408954 698614 409574 707162
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 408954 -3226 409574 14058
rect 408954 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 409574 -3226
rect 408954 -3546 409574 -3462
rect 408954 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 409574 -3546
rect 408954 -7654 409574 -3782
rect 412674 708678 413294 711590
rect 412674 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 413294 708678
rect 412674 708358 413294 708442
rect 412674 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 413294 708358
rect 412674 666334 413294 708122
rect 412674 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 413294 666334
rect 412674 666014 413294 666098
rect 412674 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 413294 666014
rect 412674 630334 413294 665778
rect 412674 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 413294 630334
rect 412674 630014 413294 630098
rect 412674 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 413294 630014
rect 412674 594334 413294 629778
rect 412674 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 413294 594334
rect 412674 594014 413294 594098
rect 412674 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 413294 594014
rect 412674 558334 413294 593778
rect 412674 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 413294 558334
rect 412674 558014 413294 558098
rect 412674 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 413294 558014
rect 412674 522334 413294 557778
rect 412674 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 413294 522334
rect 412674 522014 413294 522098
rect 412674 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 413294 522014
rect 412674 486334 413294 521778
rect 412674 486098 412706 486334
rect 412942 486098 413026 486334
rect 413262 486098 413294 486334
rect 412674 486014 413294 486098
rect 412674 485778 412706 486014
rect 412942 485778 413026 486014
rect 413262 485778 413294 486014
rect 412674 450334 413294 485778
rect 412674 450098 412706 450334
rect 412942 450098 413026 450334
rect 413262 450098 413294 450334
rect 412674 450014 413294 450098
rect 412674 449778 412706 450014
rect 412942 449778 413026 450014
rect 413262 449778 413294 450014
rect 412674 414334 413294 449778
rect 412674 414098 412706 414334
rect 412942 414098 413026 414334
rect 413262 414098 413294 414334
rect 412674 414014 413294 414098
rect 412674 413778 412706 414014
rect 412942 413778 413026 414014
rect 413262 413778 413294 414014
rect 412674 378334 413294 413778
rect 412674 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 413294 378334
rect 412674 378014 413294 378098
rect 412674 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 413294 378014
rect 412674 342334 413294 377778
rect 412674 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 413294 342334
rect 412674 342014 413294 342098
rect 412674 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 413294 342014
rect 412674 306334 413294 341778
rect 412674 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 413294 306334
rect 412674 306014 413294 306098
rect 412674 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 413294 306014
rect 412674 270334 413294 305778
rect 412674 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 413294 270334
rect 412674 270014 413294 270098
rect 412674 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 413294 270014
rect 412674 234334 413294 269778
rect 412674 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 413294 234334
rect 412674 234014 413294 234098
rect 412674 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 413294 234014
rect 412674 198334 413294 233778
rect 412674 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 413294 198334
rect 412674 198014 413294 198098
rect 412674 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 413294 198014
rect 412674 162334 413294 197778
rect 412674 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 413294 162334
rect 412674 162014 413294 162098
rect 412674 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 413294 162014
rect 412674 126334 413294 161778
rect 412674 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 413294 126334
rect 412674 126014 413294 126098
rect 412674 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 413294 126014
rect 412674 90334 413294 125778
rect 412674 90098 412706 90334
rect 412942 90098 413026 90334
rect 413262 90098 413294 90334
rect 412674 90014 413294 90098
rect 412674 89778 412706 90014
rect 412942 89778 413026 90014
rect 413262 89778 413294 90014
rect 412674 54334 413294 89778
rect 412674 54098 412706 54334
rect 412942 54098 413026 54334
rect 413262 54098 413294 54334
rect 412674 54014 413294 54098
rect 412674 53778 412706 54014
rect 412942 53778 413026 54014
rect 413262 53778 413294 54014
rect 412674 18334 413294 53778
rect 412674 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 413294 18334
rect 412674 18014 413294 18098
rect 412674 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 413294 18014
rect 412674 -4186 413294 17778
rect 412674 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 413294 -4186
rect 412674 -4506 413294 -4422
rect 412674 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 413294 -4506
rect 412674 -7654 413294 -4742
rect 416394 709638 417014 711590
rect 416394 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 417014 709638
rect 416394 709318 417014 709402
rect 416394 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 417014 709318
rect 416394 670054 417014 709082
rect 416394 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 417014 670054
rect 416394 669734 417014 669818
rect 416394 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 417014 669734
rect 416394 634054 417014 669498
rect 416394 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 417014 634054
rect 416394 633734 417014 633818
rect 416394 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 417014 633734
rect 416394 598054 417014 633498
rect 416394 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 417014 598054
rect 416394 597734 417014 597818
rect 416394 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 417014 597734
rect 416394 562054 417014 597498
rect 416394 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 417014 562054
rect 416394 561734 417014 561818
rect 416394 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 417014 561734
rect 416394 526054 417014 561498
rect 416394 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 417014 526054
rect 416394 525734 417014 525818
rect 416394 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 417014 525734
rect 416394 490054 417014 525498
rect 416394 489818 416426 490054
rect 416662 489818 416746 490054
rect 416982 489818 417014 490054
rect 416394 489734 417014 489818
rect 416394 489498 416426 489734
rect 416662 489498 416746 489734
rect 416982 489498 417014 489734
rect 416394 454054 417014 489498
rect 416394 453818 416426 454054
rect 416662 453818 416746 454054
rect 416982 453818 417014 454054
rect 416394 453734 417014 453818
rect 416394 453498 416426 453734
rect 416662 453498 416746 453734
rect 416982 453498 417014 453734
rect 416394 418054 417014 453498
rect 416394 417818 416426 418054
rect 416662 417818 416746 418054
rect 416982 417818 417014 418054
rect 416394 417734 417014 417818
rect 416394 417498 416426 417734
rect 416662 417498 416746 417734
rect 416982 417498 417014 417734
rect 416394 382054 417014 417498
rect 416394 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 417014 382054
rect 416394 381734 417014 381818
rect 416394 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 417014 381734
rect 416394 346054 417014 381498
rect 416394 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 417014 346054
rect 416394 345734 417014 345818
rect 416394 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 417014 345734
rect 416394 310054 417014 345498
rect 416394 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 417014 310054
rect 416394 309734 417014 309818
rect 416394 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 417014 309734
rect 416394 274054 417014 309498
rect 416394 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 417014 274054
rect 416394 273734 417014 273818
rect 416394 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 417014 273734
rect 416394 238054 417014 273498
rect 416394 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 417014 238054
rect 416394 237734 417014 237818
rect 416394 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 417014 237734
rect 416394 202054 417014 237498
rect 416394 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 417014 202054
rect 416394 201734 417014 201818
rect 416394 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 417014 201734
rect 416394 166054 417014 201498
rect 416394 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 417014 166054
rect 416394 165734 417014 165818
rect 416394 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 417014 165734
rect 416394 130054 417014 165498
rect 416394 129818 416426 130054
rect 416662 129818 416746 130054
rect 416982 129818 417014 130054
rect 416394 129734 417014 129818
rect 416394 129498 416426 129734
rect 416662 129498 416746 129734
rect 416982 129498 417014 129734
rect 416394 94054 417014 129498
rect 416394 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 417014 94054
rect 416394 93734 417014 93818
rect 416394 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 417014 93734
rect 416394 58054 417014 93498
rect 416394 57818 416426 58054
rect 416662 57818 416746 58054
rect 416982 57818 417014 58054
rect 416394 57734 417014 57818
rect 416394 57498 416426 57734
rect 416662 57498 416746 57734
rect 416982 57498 417014 57734
rect 416394 22054 417014 57498
rect 416394 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 417014 22054
rect 416394 21734 417014 21818
rect 416394 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 417014 21734
rect 416394 -5146 417014 21498
rect 416394 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 417014 -5146
rect 416394 -5466 417014 -5382
rect 416394 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 417014 -5466
rect 416394 -7654 417014 -5702
rect 420114 710598 420734 711590
rect 420114 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 420734 710598
rect 420114 710278 420734 710362
rect 420114 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 420734 710278
rect 420114 673774 420734 710042
rect 420114 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 420734 673774
rect 420114 673454 420734 673538
rect 420114 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 420734 673454
rect 420114 637774 420734 673218
rect 420114 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 420734 637774
rect 420114 637454 420734 637538
rect 420114 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 420734 637454
rect 420114 601774 420734 637218
rect 420114 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 420734 601774
rect 420114 601454 420734 601538
rect 420114 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 420734 601454
rect 420114 565774 420734 601218
rect 420114 565538 420146 565774
rect 420382 565538 420466 565774
rect 420702 565538 420734 565774
rect 420114 565454 420734 565538
rect 420114 565218 420146 565454
rect 420382 565218 420466 565454
rect 420702 565218 420734 565454
rect 420114 529774 420734 565218
rect 420114 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 420734 529774
rect 420114 529454 420734 529538
rect 420114 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 420734 529454
rect 420114 493774 420734 529218
rect 420114 493538 420146 493774
rect 420382 493538 420466 493774
rect 420702 493538 420734 493774
rect 420114 493454 420734 493538
rect 420114 493218 420146 493454
rect 420382 493218 420466 493454
rect 420702 493218 420734 493454
rect 420114 457774 420734 493218
rect 420114 457538 420146 457774
rect 420382 457538 420466 457774
rect 420702 457538 420734 457774
rect 420114 457454 420734 457538
rect 420114 457218 420146 457454
rect 420382 457218 420466 457454
rect 420702 457218 420734 457454
rect 420114 421774 420734 457218
rect 420114 421538 420146 421774
rect 420382 421538 420466 421774
rect 420702 421538 420734 421774
rect 420114 421454 420734 421538
rect 420114 421218 420146 421454
rect 420382 421218 420466 421454
rect 420702 421218 420734 421454
rect 420114 385774 420734 421218
rect 420114 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 420734 385774
rect 420114 385454 420734 385538
rect 420114 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 420734 385454
rect 420114 349774 420734 385218
rect 420114 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 420734 349774
rect 420114 349454 420734 349538
rect 420114 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 420734 349454
rect 420114 313774 420734 349218
rect 420114 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 420734 313774
rect 420114 313454 420734 313538
rect 420114 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 420734 313454
rect 420114 277774 420734 313218
rect 420114 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 420734 277774
rect 420114 277454 420734 277538
rect 420114 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 420734 277454
rect 420114 241774 420734 277218
rect 420114 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 420734 241774
rect 420114 241454 420734 241538
rect 420114 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 420734 241454
rect 420114 205774 420734 241218
rect 420114 205538 420146 205774
rect 420382 205538 420466 205774
rect 420702 205538 420734 205774
rect 420114 205454 420734 205538
rect 420114 205218 420146 205454
rect 420382 205218 420466 205454
rect 420702 205218 420734 205454
rect 420114 169774 420734 205218
rect 420114 169538 420146 169774
rect 420382 169538 420466 169774
rect 420702 169538 420734 169774
rect 420114 169454 420734 169538
rect 420114 169218 420146 169454
rect 420382 169218 420466 169454
rect 420702 169218 420734 169454
rect 420114 133774 420734 169218
rect 420114 133538 420146 133774
rect 420382 133538 420466 133774
rect 420702 133538 420734 133774
rect 420114 133454 420734 133538
rect 420114 133218 420146 133454
rect 420382 133218 420466 133454
rect 420702 133218 420734 133454
rect 420114 97774 420734 133218
rect 420114 97538 420146 97774
rect 420382 97538 420466 97774
rect 420702 97538 420734 97774
rect 420114 97454 420734 97538
rect 420114 97218 420146 97454
rect 420382 97218 420466 97454
rect 420702 97218 420734 97454
rect 420114 61774 420734 97218
rect 420114 61538 420146 61774
rect 420382 61538 420466 61774
rect 420702 61538 420734 61774
rect 420114 61454 420734 61538
rect 420114 61218 420146 61454
rect 420382 61218 420466 61454
rect 420702 61218 420734 61454
rect 420114 25774 420734 61218
rect 420114 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 420734 25774
rect 420114 25454 420734 25538
rect 420114 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 420734 25454
rect 420114 -6106 420734 25218
rect 420114 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 420734 -6106
rect 420114 -6426 420734 -6342
rect 420114 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 420734 -6426
rect 420114 -7654 420734 -6662
rect 423834 711558 424454 711590
rect 423834 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 424454 711558
rect 423834 711238 424454 711322
rect 423834 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 424454 711238
rect 423834 677494 424454 711002
rect 423834 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 424454 677494
rect 423834 677174 424454 677258
rect 423834 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 424454 677174
rect 423834 641494 424454 676938
rect 423834 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 424454 641494
rect 423834 641174 424454 641258
rect 423834 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 424454 641174
rect 423834 605494 424454 640938
rect 423834 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 424454 605494
rect 423834 605174 424454 605258
rect 423834 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 424454 605174
rect 423834 569494 424454 604938
rect 423834 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 424454 569494
rect 423834 569174 424454 569258
rect 423834 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 424454 569174
rect 423834 533494 424454 568938
rect 423834 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 424454 533494
rect 423834 533174 424454 533258
rect 423834 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 424454 533174
rect 423834 497494 424454 532938
rect 423834 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 424454 497494
rect 423834 497174 424454 497258
rect 423834 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 424454 497174
rect 423834 461494 424454 496938
rect 423834 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 424454 461494
rect 423834 461174 424454 461258
rect 423834 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 424454 461174
rect 423834 425494 424454 460938
rect 423834 425258 423866 425494
rect 424102 425258 424186 425494
rect 424422 425258 424454 425494
rect 423834 425174 424454 425258
rect 423834 424938 423866 425174
rect 424102 424938 424186 425174
rect 424422 424938 424454 425174
rect 423834 389494 424454 424938
rect 423834 389258 423866 389494
rect 424102 389258 424186 389494
rect 424422 389258 424454 389494
rect 423834 389174 424454 389258
rect 423834 388938 423866 389174
rect 424102 388938 424186 389174
rect 424422 388938 424454 389174
rect 423834 353494 424454 388938
rect 423834 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 424454 353494
rect 423834 353174 424454 353258
rect 423834 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 424454 353174
rect 423834 317494 424454 352938
rect 423834 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 424454 317494
rect 423834 317174 424454 317258
rect 423834 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 424454 317174
rect 423834 281494 424454 316938
rect 423834 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 424454 281494
rect 423834 281174 424454 281258
rect 423834 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 424454 281174
rect 423834 245494 424454 280938
rect 423834 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 424454 245494
rect 423834 245174 424454 245258
rect 423834 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 424454 245174
rect 423834 209494 424454 244938
rect 423834 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 424454 209494
rect 423834 209174 424454 209258
rect 423834 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 424454 209174
rect 423834 173494 424454 208938
rect 423834 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 424454 173494
rect 423834 173174 424454 173258
rect 423834 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 424454 173174
rect 423834 137494 424454 172938
rect 423834 137258 423866 137494
rect 424102 137258 424186 137494
rect 424422 137258 424454 137494
rect 423834 137174 424454 137258
rect 423834 136938 423866 137174
rect 424102 136938 424186 137174
rect 424422 136938 424454 137174
rect 423834 101494 424454 136938
rect 423834 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 424454 101494
rect 423834 101174 424454 101258
rect 423834 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 424454 101174
rect 423834 65494 424454 100938
rect 423834 65258 423866 65494
rect 424102 65258 424186 65494
rect 424422 65258 424454 65494
rect 423834 65174 424454 65258
rect 423834 64938 423866 65174
rect 424102 64938 424186 65174
rect 424422 64938 424454 65174
rect 423834 29494 424454 64938
rect 423834 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 424454 29494
rect 423834 29174 424454 29258
rect 423834 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 424454 29174
rect 423834 -7066 424454 28938
rect 423834 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 424454 -7066
rect 423834 -7386 424454 -7302
rect 423834 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 424454 -7386
rect 423834 -7654 424454 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 437514 705798 438134 711590
rect 437514 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 438134 705798
rect 437514 705478 438134 705562
rect 437514 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 438134 705478
rect 437514 691174 438134 705242
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -1306 438134 6618
rect 437514 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 438134 -1306
rect 437514 -1626 438134 -1542
rect 437514 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 438134 -1626
rect 437514 -7654 438134 -1862
rect 441234 706758 441854 711590
rect 441234 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 441854 706758
rect 441234 706438 441854 706522
rect 441234 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 441854 706438
rect 441234 694894 441854 706202
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -2266 441854 10338
rect 441234 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 441854 -2266
rect 441234 -2586 441854 -2502
rect 441234 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 441854 -2586
rect 441234 -7654 441854 -2822
rect 444954 707718 445574 711590
rect 444954 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 445574 707718
rect 444954 707398 445574 707482
rect 444954 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 445574 707398
rect 444954 698614 445574 707162
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 444954 -3226 445574 14058
rect 444954 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 445574 -3226
rect 444954 -3546 445574 -3462
rect 444954 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 445574 -3546
rect 444954 -7654 445574 -3782
rect 448674 708678 449294 711590
rect 448674 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 449294 708678
rect 448674 708358 449294 708442
rect 448674 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 449294 708358
rect 448674 666334 449294 708122
rect 448674 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 449294 666334
rect 448674 666014 449294 666098
rect 448674 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 449294 666014
rect 448674 630334 449294 665778
rect 448674 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 449294 630334
rect 448674 630014 449294 630098
rect 448674 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 449294 630014
rect 448674 594334 449294 629778
rect 448674 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 449294 594334
rect 448674 594014 449294 594098
rect 448674 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 449294 594014
rect 448674 558334 449294 593778
rect 448674 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 449294 558334
rect 448674 558014 449294 558098
rect 448674 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 449294 558014
rect 448674 522334 449294 557778
rect 448674 522098 448706 522334
rect 448942 522098 449026 522334
rect 449262 522098 449294 522334
rect 448674 522014 449294 522098
rect 448674 521778 448706 522014
rect 448942 521778 449026 522014
rect 449262 521778 449294 522014
rect 448674 486334 449294 521778
rect 448674 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 449294 486334
rect 448674 486014 449294 486098
rect 448674 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 449294 486014
rect 448674 450334 449294 485778
rect 448674 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 449294 450334
rect 448674 450014 449294 450098
rect 448674 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 449294 450014
rect 448674 414334 449294 449778
rect 448674 414098 448706 414334
rect 448942 414098 449026 414334
rect 449262 414098 449294 414334
rect 448674 414014 449294 414098
rect 448674 413778 448706 414014
rect 448942 413778 449026 414014
rect 449262 413778 449294 414014
rect 448674 378334 449294 413778
rect 448674 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 449294 378334
rect 448674 378014 449294 378098
rect 448674 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 449294 378014
rect 448674 342334 449294 377778
rect 448674 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 449294 342334
rect 448674 342014 449294 342098
rect 448674 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 449294 342014
rect 448674 306334 449294 341778
rect 448674 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 449294 306334
rect 448674 306014 449294 306098
rect 448674 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 449294 306014
rect 448674 270334 449294 305778
rect 448674 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 449294 270334
rect 448674 270014 449294 270098
rect 448674 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 449294 270014
rect 448674 234334 449294 269778
rect 448674 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 449294 234334
rect 448674 234014 449294 234098
rect 448674 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 449294 234014
rect 448674 198334 449294 233778
rect 448674 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 449294 198334
rect 448674 198014 449294 198098
rect 448674 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 449294 198014
rect 448674 162334 449294 197778
rect 448674 162098 448706 162334
rect 448942 162098 449026 162334
rect 449262 162098 449294 162334
rect 448674 162014 449294 162098
rect 448674 161778 448706 162014
rect 448942 161778 449026 162014
rect 449262 161778 449294 162014
rect 448674 126334 449294 161778
rect 448674 126098 448706 126334
rect 448942 126098 449026 126334
rect 449262 126098 449294 126334
rect 448674 126014 449294 126098
rect 448674 125778 448706 126014
rect 448942 125778 449026 126014
rect 449262 125778 449294 126014
rect 448674 90334 449294 125778
rect 448674 90098 448706 90334
rect 448942 90098 449026 90334
rect 449262 90098 449294 90334
rect 448674 90014 449294 90098
rect 448674 89778 448706 90014
rect 448942 89778 449026 90014
rect 449262 89778 449294 90014
rect 448674 54334 449294 89778
rect 448674 54098 448706 54334
rect 448942 54098 449026 54334
rect 449262 54098 449294 54334
rect 448674 54014 449294 54098
rect 448674 53778 448706 54014
rect 448942 53778 449026 54014
rect 449262 53778 449294 54014
rect 448674 18334 449294 53778
rect 448674 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 449294 18334
rect 448674 18014 449294 18098
rect 448674 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 449294 18014
rect 448674 -4186 449294 17778
rect 448674 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 449294 -4186
rect 448674 -4506 449294 -4422
rect 448674 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 449294 -4506
rect 448674 -7654 449294 -4742
rect 452394 709638 453014 711590
rect 452394 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 453014 709638
rect 452394 709318 453014 709402
rect 452394 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 453014 709318
rect 452394 670054 453014 709082
rect 452394 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 453014 670054
rect 452394 669734 453014 669818
rect 452394 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 453014 669734
rect 452394 634054 453014 669498
rect 452394 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 453014 634054
rect 452394 633734 453014 633818
rect 452394 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 453014 633734
rect 452394 598054 453014 633498
rect 452394 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 453014 598054
rect 452394 597734 453014 597818
rect 452394 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 453014 597734
rect 452394 562054 453014 597498
rect 452394 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 453014 562054
rect 452394 561734 453014 561818
rect 452394 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 453014 561734
rect 452394 526054 453014 561498
rect 452394 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 453014 526054
rect 452394 525734 453014 525818
rect 452394 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 453014 525734
rect 452394 490054 453014 525498
rect 452394 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 453014 490054
rect 452394 489734 453014 489818
rect 452394 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 453014 489734
rect 452394 454054 453014 489498
rect 452394 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 453818 453014 454054
rect 452394 453734 453014 453818
rect 452394 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 453014 453734
rect 452394 418054 453014 453498
rect 452394 417818 452426 418054
rect 452662 417818 452746 418054
rect 452982 417818 453014 418054
rect 452394 417734 453014 417818
rect 452394 417498 452426 417734
rect 452662 417498 452746 417734
rect 452982 417498 453014 417734
rect 452394 382054 453014 417498
rect 452394 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 453014 382054
rect 452394 381734 453014 381818
rect 452394 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 453014 381734
rect 452394 346054 453014 381498
rect 452394 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 453014 346054
rect 452394 345734 453014 345818
rect 452394 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 453014 345734
rect 452394 310054 453014 345498
rect 452394 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 453014 310054
rect 452394 309734 453014 309818
rect 452394 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 453014 309734
rect 452394 274054 453014 309498
rect 452394 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 453014 274054
rect 452394 273734 453014 273818
rect 452394 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 453014 273734
rect 452394 238054 453014 273498
rect 452394 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 453014 238054
rect 452394 237734 453014 237818
rect 452394 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 453014 237734
rect 452394 202054 453014 237498
rect 452394 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 453014 202054
rect 452394 201734 453014 201818
rect 452394 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 453014 201734
rect 452394 166054 453014 201498
rect 452394 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 453014 166054
rect 452394 165734 453014 165818
rect 452394 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 453014 165734
rect 452394 130054 453014 165498
rect 452394 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 453014 130054
rect 452394 129734 453014 129818
rect 452394 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 453014 129734
rect 452394 94054 453014 129498
rect 452394 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 453014 94054
rect 452394 93734 453014 93818
rect 452394 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 453014 93734
rect 452394 58054 453014 93498
rect 452394 57818 452426 58054
rect 452662 57818 452746 58054
rect 452982 57818 453014 58054
rect 452394 57734 453014 57818
rect 452394 57498 452426 57734
rect 452662 57498 452746 57734
rect 452982 57498 453014 57734
rect 452394 22054 453014 57498
rect 452394 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 453014 22054
rect 452394 21734 453014 21818
rect 452394 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 453014 21734
rect 452394 -5146 453014 21498
rect 452394 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 453014 -5146
rect 452394 -5466 453014 -5382
rect 452394 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 453014 -5466
rect 452394 -7654 453014 -5702
rect 456114 710598 456734 711590
rect 456114 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 456734 710598
rect 456114 710278 456734 710362
rect 456114 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 456734 710278
rect 456114 673774 456734 710042
rect 456114 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 456734 673774
rect 456114 673454 456734 673538
rect 456114 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 456734 673454
rect 456114 637774 456734 673218
rect 456114 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 456734 637774
rect 456114 637454 456734 637538
rect 456114 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 456734 637454
rect 456114 601774 456734 637218
rect 456114 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 456734 601774
rect 456114 601454 456734 601538
rect 456114 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 456734 601454
rect 456114 565774 456734 601218
rect 456114 565538 456146 565774
rect 456382 565538 456466 565774
rect 456702 565538 456734 565774
rect 456114 565454 456734 565538
rect 456114 565218 456146 565454
rect 456382 565218 456466 565454
rect 456702 565218 456734 565454
rect 456114 529774 456734 565218
rect 456114 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 456734 529774
rect 456114 529454 456734 529538
rect 456114 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 456734 529454
rect 456114 493774 456734 529218
rect 456114 493538 456146 493774
rect 456382 493538 456466 493774
rect 456702 493538 456734 493774
rect 456114 493454 456734 493538
rect 456114 493218 456146 493454
rect 456382 493218 456466 493454
rect 456702 493218 456734 493454
rect 456114 457774 456734 493218
rect 456114 457538 456146 457774
rect 456382 457538 456466 457774
rect 456702 457538 456734 457774
rect 456114 457454 456734 457538
rect 456114 457218 456146 457454
rect 456382 457218 456466 457454
rect 456702 457218 456734 457454
rect 456114 421774 456734 457218
rect 456114 421538 456146 421774
rect 456382 421538 456466 421774
rect 456702 421538 456734 421774
rect 456114 421454 456734 421538
rect 456114 421218 456146 421454
rect 456382 421218 456466 421454
rect 456702 421218 456734 421454
rect 456114 385774 456734 421218
rect 456114 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 456734 385774
rect 456114 385454 456734 385538
rect 456114 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 456734 385454
rect 456114 349774 456734 385218
rect 456114 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 456734 349774
rect 456114 349454 456734 349538
rect 456114 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 456734 349454
rect 456114 313774 456734 349218
rect 456114 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 456734 313774
rect 456114 313454 456734 313538
rect 456114 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 456734 313454
rect 456114 277774 456734 313218
rect 456114 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 456734 277774
rect 456114 277454 456734 277538
rect 456114 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 456734 277454
rect 456114 241774 456734 277218
rect 456114 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 456734 241774
rect 456114 241454 456734 241538
rect 456114 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 456734 241454
rect 456114 205774 456734 241218
rect 456114 205538 456146 205774
rect 456382 205538 456466 205774
rect 456702 205538 456734 205774
rect 456114 205454 456734 205538
rect 456114 205218 456146 205454
rect 456382 205218 456466 205454
rect 456702 205218 456734 205454
rect 456114 169774 456734 205218
rect 456114 169538 456146 169774
rect 456382 169538 456466 169774
rect 456702 169538 456734 169774
rect 456114 169454 456734 169538
rect 456114 169218 456146 169454
rect 456382 169218 456466 169454
rect 456702 169218 456734 169454
rect 456114 133774 456734 169218
rect 456114 133538 456146 133774
rect 456382 133538 456466 133774
rect 456702 133538 456734 133774
rect 456114 133454 456734 133538
rect 456114 133218 456146 133454
rect 456382 133218 456466 133454
rect 456702 133218 456734 133454
rect 456114 97774 456734 133218
rect 456114 97538 456146 97774
rect 456382 97538 456466 97774
rect 456702 97538 456734 97774
rect 456114 97454 456734 97538
rect 456114 97218 456146 97454
rect 456382 97218 456466 97454
rect 456702 97218 456734 97454
rect 456114 61774 456734 97218
rect 456114 61538 456146 61774
rect 456382 61538 456466 61774
rect 456702 61538 456734 61774
rect 456114 61454 456734 61538
rect 456114 61218 456146 61454
rect 456382 61218 456466 61454
rect 456702 61218 456734 61454
rect 456114 25774 456734 61218
rect 456114 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 456734 25774
rect 456114 25454 456734 25538
rect 456114 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 456734 25454
rect 456114 -6106 456734 25218
rect 456114 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 456734 -6106
rect 456114 -6426 456734 -6342
rect 456114 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 456734 -6426
rect 456114 -7654 456734 -6662
rect 459834 711558 460454 711590
rect 459834 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 460454 711558
rect 459834 711238 460454 711322
rect 459834 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 460454 711238
rect 459834 677494 460454 711002
rect 459834 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 460454 677494
rect 459834 677174 460454 677258
rect 459834 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 460454 677174
rect 459834 641494 460454 676938
rect 459834 641258 459866 641494
rect 460102 641258 460186 641494
rect 460422 641258 460454 641494
rect 459834 641174 460454 641258
rect 459834 640938 459866 641174
rect 460102 640938 460186 641174
rect 460422 640938 460454 641174
rect 459834 605494 460454 640938
rect 459834 605258 459866 605494
rect 460102 605258 460186 605494
rect 460422 605258 460454 605494
rect 459834 605174 460454 605258
rect 459834 604938 459866 605174
rect 460102 604938 460186 605174
rect 460422 604938 460454 605174
rect 459834 569494 460454 604938
rect 459834 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 460454 569494
rect 459834 569174 460454 569258
rect 459834 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 460454 569174
rect 459834 533494 460454 568938
rect 459834 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 460454 533494
rect 459834 533174 460454 533258
rect 459834 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 460454 533174
rect 459834 497494 460454 532938
rect 459834 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 460454 497494
rect 459834 497174 460454 497258
rect 459834 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 460454 497174
rect 459834 461494 460454 496938
rect 459834 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 460454 461494
rect 459834 461174 460454 461258
rect 459834 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 460454 461174
rect 459834 425494 460454 460938
rect 459834 425258 459866 425494
rect 460102 425258 460186 425494
rect 460422 425258 460454 425494
rect 459834 425174 460454 425258
rect 459834 424938 459866 425174
rect 460102 424938 460186 425174
rect 460422 424938 460454 425174
rect 459834 389494 460454 424938
rect 459834 389258 459866 389494
rect 460102 389258 460186 389494
rect 460422 389258 460454 389494
rect 459834 389174 460454 389258
rect 459834 388938 459866 389174
rect 460102 388938 460186 389174
rect 460422 388938 460454 389174
rect 459834 353494 460454 388938
rect 459834 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 460454 353494
rect 459834 353174 460454 353258
rect 459834 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 460454 353174
rect 459834 317494 460454 352938
rect 459834 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 460454 317494
rect 459834 317174 460454 317258
rect 459834 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 460454 317174
rect 459834 281494 460454 316938
rect 459834 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 460454 281494
rect 459834 281174 460454 281258
rect 459834 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 460454 281174
rect 459834 245494 460454 280938
rect 459834 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 460454 245494
rect 459834 245174 460454 245258
rect 459834 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 460454 245174
rect 459834 209494 460454 244938
rect 459834 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 460454 209494
rect 459834 209174 460454 209258
rect 459834 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 460454 209174
rect 459834 173494 460454 208938
rect 459834 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 460454 173494
rect 459834 173174 460454 173258
rect 459834 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 460454 173174
rect 459834 137494 460454 172938
rect 459834 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 460454 137494
rect 459834 137174 460454 137258
rect 459834 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 460454 137174
rect 459834 101494 460454 136938
rect 459834 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 460454 101494
rect 459834 101174 460454 101258
rect 459834 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 460454 101174
rect 459834 65494 460454 100938
rect 459834 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 460454 65494
rect 459834 65174 460454 65258
rect 459834 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 460454 65174
rect 459834 29494 460454 64938
rect 459834 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 460454 29494
rect 459834 29174 460454 29258
rect 459834 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 460454 29174
rect 459834 -7066 460454 28938
rect 459834 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 460454 -7066
rect 459834 -7386 460454 -7302
rect 459834 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 460454 -7386
rect 459834 -7654 460454 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 473514 705798 474134 711590
rect 473514 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 474134 705798
rect 473514 705478 474134 705562
rect 473514 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 474134 705478
rect 473514 691174 474134 705242
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -1306 474134 6618
rect 473514 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 474134 -1306
rect 473514 -1626 474134 -1542
rect 473514 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 474134 -1626
rect 473514 -7654 474134 -1862
rect 477234 706758 477854 711590
rect 477234 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 477854 706758
rect 477234 706438 477854 706522
rect 477234 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 477854 706438
rect 477234 694894 477854 706202
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -2266 477854 10338
rect 477234 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 477854 -2266
rect 477234 -2586 477854 -2502
rect 477234 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 477854 -2586
rect 477234 -7654 477854 -2822
rect 480954 707718 481574 711590
rect 480954 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 481574 707718
rect 480954 707398 481574 707482
rect 480954 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 481574 707398
rect 480954 698614 481574 707162
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 480954 -3226 481574 14058
rect 480954 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 481574 -3226
rect 480954 -3546 481574 -3462
rect 480954 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 481574 -3546
rect 480954 -7654 481574 -3782
rect 484674 708678 485294 711590
rect 484674 708442 484706 708678
rect 484942 708442 485026 708678
rect 485262 708442 485294 708678
rect 484674 708358 485294 708442
rect 484674 708122 484706 708358
rect 484942 708122 485026 708358
rect 485262 708122 485294 708358
rect 484674 666334 485294 708122
rect 484674 666098 484706 666334
rect 484942 666098 485026 666334
rect 485262 666098 485294 666334
rect 484674 666014 485294 666098
rect 484674 665778 484706 666014
rect 484942 665778 485026 666014
rect 485262 665778 485294 666014
rect 484674 630334 485294 665778
rect 484674 630098 484706 630334
rect 484942 630098 485026 630334
rect 485262 630098 485294 630334
rect 484674 630014 485294 630098
rect 484674 629778 484706 630014
rect 484942 629778 485026 630014
rect 485262 629778 485294 630014
rect 484674 594334 485294 629778
rect 484674 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 485294 594334
rect 484674 594014 485294 594098
rect 484674 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 485294 594014
rect 484674 558334 485294 593778
rect 484674 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 485294 558334
rect 484674 558014 485294 558098
rect 484674 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 485294 558014
rect 484674 522334 485294 557778
rect 484674 522098 484706 522334
rect 484942 522098 485026 522334
rect 485262 522098 485294 522334
rect 484674 522014 485294 522098
rect 484674 521778 484706 522014
rect 484942 521778 485026 522014
rect 485262 521778 485294 522014
rect 484674 486334 485294 521778
rect 484674 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 485294 486334
rect 484674 486014 485294 486098
rect 484674 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 485294 486014
rect 484674 450334 485294 485778
rect 484674 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 485294 450334
rect 484674 450014 485294 450098
rect 484674 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 485294 450014
rect 484674 414334 485294 449778
rect 484674 414098 484706 414334
rect 484942 414098 485026 414334
rect 485262 414098 485294 414334
rect 484674 414014 485294 414098
rect 484674 413778 484706 414014
rect 484942 413778 485026 414014
rect 485262 413778 485294 414014
rect 484674 378334 485294 413778
rect 484674 378098 484706 378334
rect 484942 378098 485026 378334
rect 485262 378098 485294 378334
rect 484674 378014 485294 378098
rect 484674 377778 484706 378014
rect 484942 377778 485026 378014
rect 485262 377778 485294 378014
rect 484674 342334 485294 377778
rect 484674 342098 484706 342334
rect 484942 342098 485026 342334
rect 485262 342098 485294 342334
rect 484674 342014 485294 342098
rect 484674 341778 484706 342014
rect 484942 341778 485026 342014
rect 485262 341778 485294 342014
rect 484674 306334 485294 341778
rect 484674 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 485294 306334
rect 484674 306014 485294 306098
rect 484674 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 485294 306014
rect 484674 270334 485294 305778
rect 484674 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 485294 270334
rect 484674 270014 485294 270098
rect 484674 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 485294 270014
rect 484674 234334 485294 269778
rect 484674 234098 484706 234334
rect 484942 234098 485026 234334
rect 485262 234098 485294 234334
rect 484674 234014 485294 234098
rect 484674 233778 484706 234014
rect 484942 233778 485026 234014
rect 485262 233778 485294 234014
rect 484674 198334 485294 233778
rect 484674 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 485294 198334
rect 484674 198014 485294 198098
rect 484674 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 485294 198014
rect 484674 162334 485294 197778
rect 484674 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 485294 162334
rect 484674 162014 485294 162098
rect 484674 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 485294 162014
rect 484674 126334 485294 161778
rect 484674 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 485294 126334
rect 484674 126014 485294 126098
rect 484674 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 485294 126014
rect 484674 90334 485294 125778
rect 484674 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 485294 90334
rect 484674 90014 485294 90098
rect 484674 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 485294 90014
rect 484674 54334 485294 89778
rect 484674 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 485294 54334
rect 484674 54014 485294 54098
rect 484674 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 485294 54014
rect 484674 18334 485294 53778
rect 484674 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 485294 18334
rect 484674 18014 485294 18098
rect 484674 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 485294 18014
rect 484674 -4186 485294 17778
rect 484674 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 485294 -4186
rect 484674 -4506 485294 -4422
rect 484674 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 485294 -4506
rect 484674 -7654 485294 -4742
rect 488394 709638 489014 711590
rect 488394 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 489014 709638
rect 488394 709318 489014 709402
rect 488394 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 489014 709318
rect 488394 670054 489014 709082
rect 488394 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 489014 670054
rect 488394 669734 489014 669818
rect 488394 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 489014 669734
rect 488394 634054 489014 669498
rect 488394 633818 488426 634054
rect 488662 633818 488746 634054
rect 488982 633818 489014 634054
rect 488394 633734 489014 633818
rect 488394 633498 488426 633734
rect 488662 633498 488746 633734
rect 488982 633498 489014 633734
rect 488394 598054 489014 633498
rect 488394 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 489014 598054
rect 488394 597734 489014 597818
rect 488394 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 489014 597734
rect 488394 562054 489014 597498
rect 488394 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 489014 562054
rect 488394 561734 489014 561818
rect 488394 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 489014 561734
rect 488394 526054 489014 561498
rect 488394 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 489014 526054
rect 488394 525734 489014 525818
rect 488394 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 489014 525734
rect 488394 490054 489014 525498
rect 488394 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 489014 490054
rect 488394 489734 489014 489818
rect 488394 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 489014 489734
rect 488394 454054 489014 489498
rect 488394 453818 488426 454054
rect 488662 453818 488746 454054
rect 488982 453818 489014 454054
rect 488394 453734 489014 453818
rect 488394 453498 488426 453734
rect 488662 453498 488746 453734
rect 488982 453498 489014 453734
rect 488394 418054 489014 453498
rect 488394 417818 488426 418054
rect 488662 417818 488746 418054
rect 488982 417818 489014 418054
rect 488394 417734 489014 417818
rect 488394 417498 488426 417734
rect 488662 417498 488746 417734
rect 488982 417498 489014 417734
rect 488394 382054 489014 417498
rect 488394 381818 488426 382054
rect 488662 381818 488746 382054
rect 488982 381818 489014 382054
rect 488394 381734 489014 381818
rect 488394 381498 488426 381734
rect 488662 381498 488746 381734
rect 488982 381498 489014 381734
rect 488394 346054 489014 381498
rect 488394 345818 488426 346054
rect 488662 345818 488746 346054
rect 488982 345818 489014 346054
rect 488394 345734 489014 345818
rect 488394 345498 488426 345734
rect 488662 345498 488746 345734
rect 488982 345498 489014 345734
rect 488394 310054 489014 345498
rect 488394 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 489014 310054
rect 488394 309734 489014 309818
rect 488394 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 489014 309734
rect 488394 274054 489014 309498
rect 488394 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 489014 274054
rect 488394 273734 489014 273818
rect 488394 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 489014 273734
rect 488394 238054 489014 273498
rect 488394 237818 488426 238054
rect 488662 237818 488746 238054
rect 488982 237818 489014 238054
rect 488394 237734 489014 237818
rect 488394 237498 488426 237734
rect 488662 237498 488746 237734
rect 488982 237498 489014 237734
rect 488394 202054 489014 237498
rect 488394 201818 488426 202054
rect 488662 201818 488746 202054
rect 488982 201818 489014 202054
rect 488394 201734 489014 201818
rect 488394 201498 488426 201734
rect 488662 201498 488746 201734
rect 488982 201498 489014 201734
rect 488394 166054 489014 201498
rect 488394 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 489014 166054
rect 488394 165734 489014 165818
rect 488394 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 489014 165734
rect 488394 130054 489014 165498
rect 488394 129818 488426 130054
rect 488662 129818 488746 130054
rect 488982 129818 489014 130054
rect 488394 129734 489014 129818
rect 488394 129498 488426 129734
rect 488662 129498 488746 129734
rect 488982 129498 489014 129734
rect 488394 94054 489014 129498
rect 488394 93818 488426 94054
rect 488662 93818 488746 94054
rect 488982 93818 489014 94054
rect 488394 93734 489014 93818
rect 488394 93498 488426 93734
rect 488662 93498 488746 93734
rect 488982 93498 489014 93734
rect 488394 58054 489014 93498
rect 488394 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 489014 58054
rect 488394 57734 489014 57818
rect 488394 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 489014 57734
rect 488394 22054 489014 57498
rect 488394 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 489014 22054
rect 488394 21734 489014 21818
rect 488394 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 489014 21734
rect 488394 -5146 489014 21498
rect 488394 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 489014 -5146
rect 488394 -5466 489014 -5382
rect 488394 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 489014 -5466
rect 488394 -7654 489014 -5702
rect 492114 710598 492734 711590
rect 492114 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 492734 710598
rect 492114 710278 492734 710362
rect 492114 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 492734 710278
rect 492114 673774 492734 710042
rect 492114 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 492734 673774
rect 492114 673454 492734 673538
rect 492114 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 492734 673454
rect 492114 637774 492734 673218
rect 492114 637538 492146 637774
rect 492382 637538 492466 637774
rect 492702 637538 492734 637774
rect 492114 637454 492734 637538
rect 492114 637218 492146 637454
rect 492382 637218 492466 637454
rect 492702 637218 492734 637454
rect 492114 601774 492734 637218
rect 492114 601538 492146 601774
rect 492382 601538 492466 601774
rect 492702 601538 492734 601774
rect 492114 601454 492734 601538
rect 492114 601218 492146 601454
rect 492382 601218 492466 601454
rect 492702 601218 492734 601454
rect 492114 565774 492734 601218
rect 492114 565538 492146 565774
rect 492382 565538 492466 565774
rect 492702 565538 492734 565774
rect 492114 565454 492734 565538
rect 492114 565218 492146 565454
rect 492382 565218 492466 565454
rect 492702 565218 492734 565454
rect 492114 529774 492734 565218
rect 492114 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 492734 529774
rect 492114 529454 492734 529538
rect 492114 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 492734 529454
rect 492114 493774 492734 529218
rect 492114 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 492734 493774
rect 492114 493454 492734 493538
rect 492114 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 492734 493454
rect 492114 457774 492734 493218
rect 492114 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 492734 457774
rect 492114 457454 492734 457538
rect 492114 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 492734 457454
rect 492114 421774 492734 457218
rect 492114 421538 492146 421774
rect 492382 421538 492466 421774
rect 492702 421538 492734 421774
rect 492114 421454 492734 421538
rect 492114 421218 492146 421454
rect 492382 421218 492466 421454
rect 492702 421218 492734 421454
rect 492114 385774 492734 421218
rect 492114 385538 492146 385774
rect 492382 385538 492466 385774
rect 492702 385538 492734 385774
rect 492114 385454 492734 385538
rect 492114 385218 492146 385454
rect 492382 385218 492466 385454
rect 492702 385218 492734 385454
rect 492114 349774 492734 385218
rect 492114 349538 492146 349774
rect 492382 349538 492466 349774
rect 492702 349538 492734 349774
rect 492114 349454 492734 349538
rect 492114 349218 492146 349454
rect 492382 349218 492466 349454
rect 492702 349218 492734 349454
rect 492114 313774 492734 349218
rect 492114 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 492734 313774
rect 492114 313454 492734 313538
rect 492114 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 492734 313454
rect 492114 277774 492734 313218
rect 492114 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 492734 277774
rect 492114 277454 492734 277538
rect 492114 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 492734 277454
rect 492114 241774 492734 277218
rect 492114 241538 492146 241774
rect 492382 241538 492466 241774
rect 492702 241538 492734 241774
rect 492114 241454 492734 241538
rect 492114 241218 492146 241454
rect 492382 241218 492466 241454
rect 492702 241218 492734 241454
rect 492114 205774 492734 241218
rect 492114 205538 492146 205774
rect 492382 205538 492466 205774
rect 492702 205538 492734 205774
rect 492114 205454 492734 205538
rect 492114 205218 492146 205454
rect 492382 205218 492466 205454
rect 492702 205218 492734 205454
rect 492114 169774 492734 205218
rect 492114 169538 492146 169774
rect 492382 169538 492466 169774
rect 492702 169538 492734 169774
rect 492114 169454 492734 169538
rect 492114 169218 492146 169454
rect 492382 169218 492466 169454
rect 492702 169218 492734 169454
rect 492114 133774 492734 169218
rect 492114 133538 492146 133774
rect 492382 133538 492466 133774
rect 492702 133538 492734 133774
rect 492114 133454 492734 133538
rect 492114 133218 492146 133454
rect 492382 133218 492466 133454
rect 492702 133218 492734 133454
rect 492114 97774 492734 133218
rect 492114 97538 492146 97774
rect 492382 97538 492466 97774
rect 492702 97538 492734 97774
rect 492114 97454 492734 97538
rect 492114 97218 492146 97454
rect 492382 97218 492466 97454
rect 492702 97218 492734 97454
rect 492114 61774 492734 97218
rect 492114 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 492734 61774
rect 492114 61454 492734 61538
rect 492114 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 492734 61454
rect 492114 25774 492734 61218
rect 492114 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 492734 25774
rect 492114 25454 492734 25538
rect 492114 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 492734 25454
rect 492114 -6106 492734 25218
rect 492114 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 492734 -6106
rect 492114 -6426 492734 -6342
rect 492114 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 492734 -6426
rect 492114 -7654 492734 -6662
rect 495834 711558 496454 711590
rect 495834 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 496454 711558
rect 495834 711238 496454 711322
rect 495834 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 496454 711238
rect 495834 677494 496454 711002
rect 495834 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 496454 677494
rect 495834 677174 496454 677258
rect 495834 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 496454 677174
rect 495834 641494 496454 676938
rect 495834 641258 495866 641494
rect 496102 641258 496186 641494
rect 496422 641258 496454 641494
rect 495834 641174 496454 641258
rect 495834 640938 495866 641174
rect 496102 640938 496186 641174
rect 496422 640938 496454 641174
rect 495834 605494 496454 640938
rect 495834 605258 495866 605494
rect 496102 605258 496186 605494
rect 496422 605258 496454 605494
rect 495834 605174 496454 605258
rect 495834 604938 495866 605174
rect 496102 604938 496186 605174
rect 496422 604938 496454 605174
rect 495834 569494 496454 604938
rect 495834 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 496454 569494
rect 495834 569174 496454 569258
rect 495834 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 496454 569174
rect 495834 533494 496454 568938
rect 495834 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 496454 533494
rect 495834 533174 496454 533258
rect 495834 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 496454 533174
rect 495834 497494 496454 532938
rect 495834 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 496454 497494
rect 495834 497174 496454 497258
rect 495834 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 496454 497174
rect 495834 461494 496454 496938
rect 495834 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 496454 461494
rect 495834 461174 496454 461258
rect 495834 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 496454 461174
rect 495834 425494 496454 460938
rect 495834 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 496454 425494
rect 495834 425174 496454 425258
rect 495834 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 496454 425174
rect 495834 389494 496454 424938
rect 495834 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 496454 389494
rect 495834 389174 496454 389258
rect 495834 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 496454 389174
rect 495834 353494 496454 388938
rect 495834 353258 495866 353494
rect 496102 353258 496186 353494
rect 496422 353258 496454 353494
rect 495834 353174 496454 353258
rect 495834 352938 495866 353174
rect 496102 352938 496186 353174
rect 496422 352938 496454 353174
rect 495834 317494 496454 352938
rect 495834 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 496454 317494
rect 495834 317174 496454 317258
rect 495834 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 496454 317174
rect 495834 281494 496454 316938
rect 495834 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 496454 281494
rect 495834 281174 496454 281258
rect 495834 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 496454 281174
rect 495834 245494 496454 280938
rect 495834 245258 495866 245494
rect 496102 245258 496186 245494
rect 496422 245258 496454 245494
rect 495834 245174 496454 245258
rect 495834 244938 495866 245174
rect 496102 244938 496186 245174
rect 496422 244938 496454 245174
rect 495834 209494 496454 244938
rect 495834 209258 495866 209494
rect 496102 209258 496186 209494
rect 496422 209258 496454 209494
rect 495834 209174 496454 209258
rect 495834 208938 495866 209174
rect 496102 208938 496186 209174
rect 496422 208938 496454 209174
rect 495834 173494 496454 208938
rect 495834 173258 495866 173494
rect 496102 173258 496186 173494
rect 496422 173258 496454 173494
rect 495834 173174 496454 173258
rect 495834 172938 495866 173174
rect 496102 172938 496186 173174
rect 496422 172938 496454 173174
rect 495834 137494 496454 172938
rect 495834 137258 495866 137494
rect 496102 137258 496186 137494
rect 496422 137258 496454 137494
rect 495834 137174 496454 137258
rect 495834 136938 495866 137174
rect 496102 136938 496186 137174
rect 496422 136938 496454 137174
rect 495834 101494 496454 136938
rect 495834 101258 495866 101494
rect 496102 101258 496186 101494
rect 496422 101258 496454 101494
rect 495834 101174 496454 101258
rect 495834 100938 495866 101174
rect 496102 100938 496186 101174
rect 496422 100938 496454 101174
rect 495834 65494 496454 100938
rect 495834 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 496454 65494
rect 495834 65174 496454 65258
rect 495834 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 496454 65174
rect 495834 29494 496454 64938
rect 495834 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 496454 29494
rect 495834 29174 496454 29258
rect 495834 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 496454 29174
rect 495834 -7066 496454 28938
rect 495834 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 496454 -7066
rect 495834 -7386 496454 -7302
rect 495834 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 496454 -7386
rect 495834 -7654 496454 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 509514 705798 510134 711590
rect 509514 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 510134 705798
rect 509514 705478 510134 705562
rect 509514 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 510134 705478
rect 509514 691174 510134 705242
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -1306 510134 6618
rect 509514 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 510134 -1306
rect 509514 -1626 510134 -1542
rect 509514 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 510134 -1626
rect 509514 -7654 510134 -1862
rect 513234 706758 513854 711590
rect 513234 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 513854 706758
rect 513234 706438 513854 706522
rect 513234 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 513854 706438
rect 513234 694894 513854 706202
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -2266 513854 10338
rect 513234 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 513854 -2266
rect 513234 -2586 513854 -2502
rect 513234 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 513854 -2586
rect 513234 -7654 513854 -2822
rect 516954 707718 517574 711590
rect 516954 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 517574 707718
rect 516954 707398 517574 707482
rect 516954 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 517574 707398
rect 516954 698614 517574 707162
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 516954 -3226 517574 14058
rect 516954 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 517574 -3226
rect 516954 -3546 517574 -3462
rect 516954 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 517574 -3546
rect 516954 -7654 517574 -3782
rect 520674 708678 521294 711590
rect 520674 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 521294 708678
rect 520674 708358 521294 708442
rect 520674 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 521294 708358
rect 520674 666334 521294 708122
rect 520674 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 521294 666334
rect 520674 666014 521294 666098
rect 520674 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 521294 666014
rect 520674 630334 521294 665778
rect 520674 630098 520706 630334
rect 520942 630098 521026 630334
rect 521262 630098 521294 630334
rect 520674 630014 521294 630098
rect 520674 629778 520706 630014
rect 520942 629778 521026 630014
rect 521262 629778 521294 630014
rect 520674 594334 521294 629778
rect 520674 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 521294 594334
rect 520674 594014 521294 594098
rect 520674 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 521294 594014
rect 520674 558334 521294 593778
rect 520674 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 521294 558334
rect 520674 558014 521294 558098
rect 520674 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 521294 558014
rect 520674 522334 521294 557778
rect 520674 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 521294 522334
rect 520674 522014 521294 522098
rect 520674 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 521294 522014
rect 520674 486334 521294 521778
rect 520674 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 521294 486334
rect 520674 486014 521294 486098
rect 520674 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 521294 486014
rect 520674 450334 521294 485778
rect 520674 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 521294 450334
rect 520674 450014 521294 450098
rect 520674 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 521294 450014
rect 520674 414334 521294 449778
rect 520674 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 521294 414334
rect 520674 414014 521294 414098
rect 520674 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 521294 414014
rect 520674 378334 521294 413778
rect 520674 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378098 521294 378334
rect 520674 378014 521294 378098
rect 520674 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 377778 521294 378014
rect 520674 342334 521294 377778
rect 520674 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 521294 342334
rect 520674 342014 521294 342098
rect 520674 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 521294 342014
rect 520674 306334 521294 341778
rect 520674 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 521294 306334
rect 520674 306014 521294 306098
rect 520674 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 521294 306014
rect 520674 270334 521294 305778
rect 520674 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 521294 270334
rect 520674 270014 521294 270098
rect 520674 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 521294 270014
rect 520674 234334 521294 269778
rect 520674 234098 520706 234334
rect 520942 234098 521026 234334
rect 521262 234098 521294 234334
rect 520674 234014 521294 234098
rect 520674 233778 520706 234014
rect 520942 233778 521026 234014
rect 521262 233778 521294 234014
rect 520674 198334 521294 233778
rect 520674 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 521294 198334
rect 520674 198014 521294 198098
rect 520674 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 521294 198014
rect 520674 162334 521294 197778
rect 520674 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 521294 162334
rect 520674 162014 521294 162098
rect 520674 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 521294 162014
rect 520674 126334 521294 161778
rect 520674 126098 520706 126334
rect 520942 126098 521026 126334
rect 521262 126098 521294 126334
rect 520674 126014 521294 126098
rect 520674 125778 520706 126014
rect 520942 125778 521026 126014
rect 521262 125778 521294 126014
rect 520674 90334 521294 125778
rect 520674 90098 520706 90334
rect 520942 90098 521026 90334
rect 521262 90098 521294 90334
rect 520674 90014 521294 90098
rect 520674 89778 520706 90014
rect 520942 89778 521026 90014
rect 521262 89778 521294 90014
rect 520674 54334 521294 89778
rect 520674 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 521294 54334
rect 520674 54014 521294 54098
rect 520674 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 521294 54014
rect 520674 18334 521294 53778
rect 520674 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 521294 18334
rect 520674 18014 521294 18098
rect 520674 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 521294 18014
rect 520674 -4186 521294 17778
rect 520674 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 521294 -4186
rect 520674 -4506 521294 -4422
rect 520674 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 521294 -4506
rect 520674 -7654 521294 -4742
rect 524394 709638 525014 711590
rect 524394 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 525014 709638
rect 524394 709318 525014 709402
rect 524394 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 525014 709318
rect 524394 670054 525014 709082
rect 524394 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 525014 670054
rect 524394 669734 525014 669818
rect 524394 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 525014 669734
rect 524394 634054 525014 669498
rect 524394 633818 524426 634054
rect 524662 633818 524746 634054
rect 524982 633818 525014 634054
rect 524394 633734 525014 633818
rect 524394 633498 524426 633734
rect 524662 633498 524746 633734
rect 524982 633498 525014 633734
rect 524394 598054 525014 633498
rect 524394 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 525014 598054
rect 524394 597734 525014 597818
rect 524394 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 525014 597734
rect 524394 562054 525014 597498
rect 524394 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 525014 562054
rect 524394 561734 525014 561818
rect 524394 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 525014 561734
rect 524394 526054 525014 561498
rect 524394 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 525014 526054
rect 524394 525734 525014 525818
rect 524394 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 525014 525734
rect 524394 490054 525014 525498
rect 524394 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 525014 490054
rect 524394 489734 525014 489818
rect 524394 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 525014 489734
rect 524394 454054 525014 489498
rect 524394 453818 524426 454054
rect 524662 453818 524746 454054
rect 524982 453818 525014 454054
rect 524394 453734 525014 453818
rect 524394 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 525014 453734
rect 524394 418054 525014 453498
rect 524394 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 525014 418054
rect 524394 417734 525014 417818
rect 524394 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 525014 417734
rect 524394 382054 525014 417498
rect 524394 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 525014 382054
rect 524394 381734 525014 381818
rect 524394 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 525014 381734
rect 524394 346054 525014 381498
rect 524394 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 525014 346054
rect 524394 345734 525014 345818
rect 524394 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 525014 345734
rect 524394 310054 525014 345498
rect 524394 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 525014 310054
rect 524394 309734 525014 309818
rect 524394 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 525014 309734
rect 524394 274054 525014 309498
rect 524394 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 525014 274054
rect 524394 273734 525014 273818
rect 524394 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 525014 273734
rect 524394 238054 525014 273498
rect 524394 237818 524426 238054
rect 524662 237818 524746 238054
rect 524982 237818 525014 238054
rect 524394 237734 525014 237818
rect 524394 237498 524426 237734
rect 524662 237498 524746 237734
rect 524982 237498 525014 237734
rect 524394 202054 525014 237498
rect 524394 201818 524426 202054
rect 524662 201818 524746 202054
rect 524982 201818 525014 202054
rect 524394 201734 525014 201818
rect 524394 201498 524426 201734
rect 524662 201498 524746 201734
rect 524982 201498 525014 201734
rect 524394 166054 525014 201498
rect 524394 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 525014 166054
rect 524394 165734 525014 165818
rect 524394 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 525014 165734
rect 524394 130054 525014 165498
rect 524394 129818 524426 130054
rect 524662 129818 524746 130054
rect 524982 129818 525014 130054
rect 524394 129734 525014 129818
rect 524394 129498 524426 129734
rect 524662 129498 524746 129734
rect 524982 129498 525014 129734
rect 524394 94054 525014 129498
rect 524394 93818 524426 94054
rect 524662 93818 524746 94054
rect 524982 93818 525014 94054
rect 524394 93734 525014 93818
rect 524394 93498 524426 93734
rect 524662 93498 524746 93734
rect 524982 93498 525014 93734
rect 524394 58054 525014 93498
rect 524394 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 525014 58054
rect 524394 57734 525014 57818
rect 524394 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 525014 57734
rect 524394 22054 525014 57498
rect 524394 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 525014 22054
rect 524394 21734 525014 21818
rect 524394 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 525014 21734
rect 524394 -5146 525014 21498
rect 524394 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 525014 -5146
rect 524394 -5466 525014 -5382
rect 524394 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 525014 -5466
rect 524394 -7654 525014 -5702
rect 528114 710598 528734 711590
rect 528114 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 528734 710598
rect 528114 710278 528734 710362
rect 528114 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 528734 710278
rect 528114 673774 528734 710042
rect 528114 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 528734 673774
rect 528114 673454 528734 673538
rect 528114 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 528734 673454
rect 528114 637774 528734 673218
rect 528114 637538 528146 637774
rect 528382 637538 528466 637774
rect 528702 637538 528734 637774
rect 528114 637454 528734 637538
rect 528114 637218 528146 637454
rect 528382 637218 528466 637454
rect 528702 637218 528734 637454
rect 528114 601774 528734 637218
rect 528114 601538 528146 601774
rect 528382 601538 528466 601774
rect 528702 601538 528734 601774
rect 528114 601454 528734 601538
rect 528114 601218 528146 601454
rect 528382 601218 528466 601454
rect 528702 601218 528734 601454
rect 528114 565774 528734 601218
rect 528114 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 528734 565774
rect 528114 565454 528734 565538
rect 528114 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 528734 565454
rect 528114 529774 528734 565218
rect 528114 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 528734 529774
rect 528114 529454 528734 529538
rect 528114 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 528734 529454
rect 528114 493774 528734 529218
rect 528114 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 528734 493774
rect 528114 493454 528734 493538
rect 528114 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 528734 493454
rect 528114 457774 528734 493218
rect 528114 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 528734 457774
rect 528114 457454 528734 457538
rect 528114 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 528734 457454
rect 528114 421774 528734 457218
rect 528114 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 528734 421774
rect 528114 421454 528734 421538
rect 528114 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 528734 421454
rect 528114 385774 528734 421218
rect 528114 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 528734 385774
rect 528114 385454 528734 385538
rect 528114 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 528734 385454
rect 528114 349774 528734 385218
rect 528114 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 528734 349774
rect 528114 349454 528734 349538
rect 528114 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 528734 349454
rect 528114 313774 528734 349218
rect 528114 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 528734 313774
rect 528114 313454 528734 313538
rect 528114 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 528734 313454
rect 528114 277774 528734 313218
rect 528114 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 528734 277774
rect 528114 277454 528734 277538
rect 528114 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 528734 277454
rect 528114 241774 528734 277218
rect 528114 241538 528146 241774
rect 528382 241538 528466 241774
rect 528702 241538 528734 241774
rect 528114 241454 528734 241538
rect 528114 241218 528146 241454
rect 528382 241218 528466 241454
rect 528702 241218 528734 241454
rect 528114 205774 528734 241218
rect 528114 205538 528146 205774
rect 528382 205538 528466 205774
rect 528702 205538 528734 205774
rect 528114 205454 528734 205538
rect 528114 205218 528146 205454
rect 528382 205218 528466 205454
rect 528702 205218 528734 205454
rect 528114 169774 528734 205218
rect 528114 169538 528146 169774
rect 528382 169538 528466 169774
rect 528702 169538 528734 169774
rect 528114 169454 528734 169538
rect 528114 169218 528146 169454
rect 528382 169218 528466 169454
rect 528702 169218 528734 169454
rect 528114 133774 528734 169218
rect 528114 133538 528146 133774
rect 528382 133538 528466 133774
rect 528702 133538 528734 133774
rect 528114 133454 528734 133538
rect 528114 133218 528146 133454
rect 528382 133218 528466 133454
rect 528702 133218 528734 133454
rect 528114 97774 528734 133218
rect 528114 97538 528146 97774
rect 528382 97538 528466 97774
rect 528702 97538 528734 97774
rect 528114 97454 528734 97538
rect 528114 97218 528146 97454
rect 528382 97218 528466 97454
rect 528702 97218 528734 97454
rect 528114 61774 528734 97218
rect 528114 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 528734 61774
rect 528114 61454 528734 61538
rect 528114 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 528734 61454
rect 528114 25774 528734 61218
rect 528114 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 528734 25774
rect 528114 25454 528734 25538
rect 528114 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 528734 25454
rect 528114 -6106 528734 25218
rect 528114 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 528734 -6106
rect 528114 -6426 528734 -6342
rect 528114 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 528734 -6426
rect 528114 -7654 528734 -6662
rect 531834 711558 532454 711590
rect 531834 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 532454 711558
rect 531834 711238 532454 711322
rect 531834 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 532454 711238
rect 531834 677494 532454 711002
rect 531834 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 532454 677494
rect 531834 677174 532454 677258
rect 531834 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 532454 677174
rect 531834 641494 532454 676938
rect 531834 641258 531866 641494
rect 532102 641258 532186 641494
rect 532422 641258 532454 641494
rect 531834 641174 532454 641258
rect 531834 640938 531866 641174
rect 532102 640938 532186 641174
rect 532422 640938 532454 641174
rect 531834 605494 532454 640938
rect 531834 605258 531866 605494
rect 532102 605258 532186 605494
rect 532422 605258 532454 605494
rect 531834 605174 532454 605258
rect 531834 604938 531866 605174
rect 532102 604938 532186 605174
rect 532422 604938 532454 605174
rect 531834 569494 532454 604938
rect 531834 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 532454 569494
rect 531834 569174 532454 569258
rect 531834 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 532454 569174
rect 531834 533494 532454 568938
rect 531834 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 532454 533494
rect 531834 533174 532454 533258
rect 531834 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 532454 533174
rect 531834 497494 532454 532938
rect 531834 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 532454 497494
rect 531834 497174 532454 497258
rect 531834 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 532454 497174
rect 531834 461494 532454 496938
rect 531834 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 532454 461494
rect 531834 461174 532454 461258
rect 531834 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 532454 461174
rect 531834 425494 532454 460938
rect 531834 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 532454 425494
rect 531834 425174 532454 425258
rect 531834 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 532454 425174
rect 531834 389494 532454 424938
rect 531834 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 532454 389494
rect 531834 389174 532454 389258
rect 531834 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 532454 389174
rect 531834 353494 532454 388938
rect 531834 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 532454 353494
rect 531834 353174 532454 353258
rect 531834 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 532454 353174
rect 531834 317494 532454 352938
rect 531834 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 532454 317494
rect 531834 317174 532454 317258
rect 531834 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 532454 317174
rect 531834 281494 532454 316938
rect 531834 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 532454 281494
rect 531834 281174 532454 281258
rect 531834 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 532454 281174
rect 531834 245494 532454 280938
rect 531834 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 532454 245494
rect 531834 245174 532454 245258
rect 531834 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 532454 245174
rect 531834 209494 532454 244938
rect 531834 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 532454 209494
rect 531834 209174 532454 209258
rect 531834 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 532454 209174
rect 531834 173494 532454 208938
rect 531834 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 532454 173494
rect 531834 173174 532454 173258
rect 531834 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 532454 173174
rect 531834 137494 532454 172938
rect 531834 137258 531866 137494
rect 532102 137258 532186 137494
rect 532422 137258 532454 137494
rect 531834 137174 532454 137258
rect 531834 136938 531866 137174
rect 532102 136938 532186 137174
rect 532422 136938 532454 137174
rect 531834 101494 532454 136938
rect 531834 101258 531866 101494
rect 532102 101258 532186 101494
rect 532422 101258 532454 101494
rect 531834 101174 532454 101258
rect 531834 100938 531866 101174
rect 532102 100938 532186 101174
rect 532422 100938 532454 101174
rect 531834 65494 532454 100938
rect 531834 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 532454 65494
rect 531834 65174 532454 65258
rect 531834 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 532454 65174
rect 531834 29494 532454 64938
rect 531834 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 532454 29494
rect 531834 29174 532454 29258
rect 531834 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 532454 29174
rect 531834 -7066 532454 28938
rect 531834 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 532454 -7066
rect 531834 -7386 532454 -7302
rect 531834 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 532454 -7386
rect 531834 -7654 532454 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 545514 705798 546134 711590
rect 545514 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 546134 705798
rect 545514 705478 546134 705562
rect 545514 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 546134 705478
rect 545514 691174 546134 705242
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -1306 546134 6618
rect 545514 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 546134 -1306
rect 545514 -1626 546134 -1542
rect 545514 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 546134 -1626
rect 545514 -7654 546134 -1862
rect 549234 706758 549854 711590
rect 549234 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 549854 706758
rect 549234 706438 549854 706522
rect 549234 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 549854 706438
rect 549234 694894 549854 706202
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -2266 549854 10338
rect 549234 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 549854 -2266
rect 549234 -2586 549854 -2502
rect 549234 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 549854 -2586
rect 549234 -7654 549854 -2822
rect 552954 707718 553574 711590
rect 552954 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 553574 707718
rect 552954 707398 553574 707482
rect 552954 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 553574 707398
rect 552954 698614 553574 707162
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 552954 -3226 553574 14058
rect 552954 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 553574 -3226
rect 552954 -3546 553574 -3462
rect 552954 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 553574 -3546
rect 552954 -7654 553574 -3782
rect 556674 708678 557294 711590
rect 556674 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 557294 708678
rect 556674 708358 557294 708442
rect 556674 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 557294 708358
rect 556674 666334 557294 708122
rect 556674 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 557294 666334
rect 556674 666014 557294 666098
rect 556674 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 557294 666014
rect 556674 630334 557294 665778
rect 556674 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 557294 630334
rect 556674 630014 557294 630098
rect 556674 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 557294 630014
rect 556674 594334 557294 629778
rect 556674 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 557294 594334
rect 556674 594014 557294 594098
rect 556674 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 557294 594014
rect 556674 558334 557294 593778
rect 556674 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 557294 558334
rect 556674 558014 557294 558098
rect 556674 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 557294 558014
rect 556674 522334 557294 557778
rect 556674 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 557294 522334
rect 556674 522014 557294 522098
rect 556674 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 557294 522014
rect 556674 486334 557294 521778
rect 556674 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 557294 486334
rect 556674 486014 557294 486098
rect 556674 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 557294 486014
rect 556674 450334 557294 485778
rect 556674 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 557294 450334
rect 556674 450014 557294 450098
rect 556674 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 557294 450014
rect 556674 414334 557294 449778
rect 556674 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 557294 414334
rect 556674 414014 557294 414098
rect 556674 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 557294 414014
rect 556674 378334 557294 413778
rect 556674 378098 556706 378334
rect 556942 378098 557026 378334
rect 557262 378098 557294 378334
rect 556674 378014 557294 378098
rect 556674 377778 556706 378014
rect 556942 377778 557026 378014
rect 557262 377778 557294 378014
rect 556674 342334 557294 377778
rect 556674 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 557294 342334
rect 556674 342014 557294 342098
rect 556674 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 557294 342014
rect 556674 306334 557294 341778
rect 556674 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 557294 306334
rect 556674 306014 557294 306098
rect 556674 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 557294 306014
rect 556674 270334 557294 305778
rect 556674 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 557294 270334
rect 556674 270014 557294 270098
rect 556674 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 557294 270014
rect 556674 234334 557294 269778
rect 556674 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 557294 234334
rect 556674 234014 557294 234098
rect 556674 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 557294 234014
rect 556674 198334 557294 233778
rect 556674 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 557294 198334
rect 556674 198014 557294 198098
rect 556674 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 557294 198014
rect 556674 162334 557294 197778
rect 556674 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 557294 162334
rect 556674 162014 557294 162098
rect 556674 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 557294 162014
rect 556674 126334 557294 161778
rect 556674 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 557294 126334
rect 556674 126014 557294 126098
rect 556674 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 557294 126014
rect 556674 90334 557294 125778
rect 556674 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 557294 90334
rect 556674 90014 557294 90098
rect 556674 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 557294 90014
rect 556674 54334 557294 89778
rect 556674 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 557294 54334
rect 556674 54014 557294 54098
rect 556674 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 557294 54014
rect 556674 18334 557294 53778
rect 556674 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 557294 18334
rect 556674 18014 557294 18098
rect 556674 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 557294 18014
rect 556674 -4186 557294 17778
rect 556674 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 557294 -4186
rect 556674 -4506 557294 -4422
rect 556674 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 557294 -4506
rect 556674 -7654 557294 -4742
rect 560394 709638 561014 711590
rect 560394 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 561014 709638
rect 560394 709318 561014 709402
rect 560394 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 561014 709318
rect 560394 670054 561014 709082
rect 560394 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 561014 670054
rect 560394 669734 561014 669818
rect 560394 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 561014 669734
rect 560394 634054 561014 669498
rect 560394 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 561014 634054
rect 560394 633734 561014 633818
rect 560394 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 561014 633734
rect 560394 598054 561014 633498
rect 560394 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 561014 598054
rect 560394 597734 561014 597818
rect 560394 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 561014 597734
rect 560394 562054 561014 597498
rect 560394 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 561014 562054
rect 560394 561734 561014 561818
rect 560394 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 561014 561734
rect 560394 526054 561014 561498
rect 560394 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 561014 526054
rect 560394 525734 561014 525818
rect 560394 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 561014 525734
rect 560394 490054 561014 525498
rect 560394 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 561014 490054
rect 560394 489734 561014 489818
rect 560394 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 561014 489734
rect 560394 454054 561014 489498
rect 560394 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 561014 454054
rect 560394 453734 561014 453818
rect 560394 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 561014 453734
rect 560394 418054 561014 453498
rect 560394 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 561014 418054
rect 560394 417734 561014 417818
rect 560394 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 561014 417734
rect 560394 382054 561014 417498
rect 560394 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 561014 382054
rect 560394 381734 561014 381818
rect 560394 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 561014 381734
rect 560394 346054 561014 381498
rect 560394 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 561014 346054
rect 560394 345734 561014 345818
rect 560394 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 561014 345734
rect 560394 310054 561014 345498
rect 560394 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 561014 310054
rect 560394 309734 561014 309818
rect 560394 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 561014 309734
rect 560394 274054 561014 309498
rect 560394 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 561014 274054
rect 560394 273734 561014 273818
rect 560394 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 561014 273734
rect 560394 238054 561014 273498
rect 560394 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 561014 238054
rect 560394 237734 561014 237818
rect 560394 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 561014 237734
rect 560394 202054 561014 237498
rect 560394 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 561014 202054
rect 560394 201734 561014 201818
rect 560394 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 561014 201734
rect 560394 166054 561014 201498
rect 560394 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 561014 166054
rect 560394 165734 561014 165818
rect 560394 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 561014 165734
rect 560394 130054 561014 165498
rect 560394 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 561014 130054
rect 560394 129734 561014 129818
rect 560394 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 561014 129734
rect 560394 94054 561014 129498
rect 560394 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 561014 94054
rect 560394 93734 561014 93818
rect 560394 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 561014 93734
rect 560394 58054 561014 93498
rect 560394 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 561014 58054
rect 560394 57734 561014 57818
rect 560394 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 561014 57734
rect 560394 22054 561014 57498
rect 560394 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 561014 22054
rect 560394 21734 561014 21818
rect 560394 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 561014 21734
rect 560394 -5146 561014 21498
rect 560394 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 561014 -5146
rect 560394 -5466 561014 -5382
rect 560394 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 561014 -5466
rect 560394 -7654 561014 -5702
rect 564114 710598 564734 711590
rect 564114 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 564734 710598
rect 564114 710278 564734 710362
rect 564114 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 564734 710278
rect 564114 673774 564734 710042
rect 564114 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 564734 673774
rect 564114 673454 564734 673538
rect 564114 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 564734 673454
rect 564114 637774 564734 673218
rect 564114 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 564734 637774
rect 564114 637454 564734 637538
rect 564114 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 564734 637454
rect 564114 601774 564734 637218
rect 564114 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 564734 601774
rect 564114 601454 564734 601538
rect 564114 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 564734 601454
rect 564114 565774 564734 601218
rect 564114 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 564734 565774
rect 564114 565454 564734 565538
rect 564114 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 564734 565454
rect 564114 529774 564734 565218
rect 564114 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 564734 529774
rect 564114 529454 564734 529538
rect 564114 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 564734 529454
rect 564114 493774 564734 529218
rect 564114 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 564734 493774
rect 564114 493454 564734 493538
rect 564114 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 564734 493454
rect 564114 457774 564734 493218
rect 564114 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 564734 457774
rect 564114 457454 564734 457538
rect 564114 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 564734 457454
rect 564114 421774 564734 457218
rect 564114 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 564734 421774
rect 564114 421454 564734 421538
rect 564114 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 564734 421454
rect 564114 385774 564734 421218
rect 564114 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 564734 385774
rect 564114 385454 564734 385538
rect 564114 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 564734 385454
rect 564114 349774 564734 385218
rect 564114 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 564734 349774
rect 564114 349454 564734 349538
rect 564114 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 564734 349454
rect 564114 313774 564734 349218
rect 564114 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 564734 313774
rect 564114 313454 564734 313538
rect 564114 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 564734 313454
rect 564114 277774 564734 313218
rect 564114 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 564734 277774
rect 564114 277454 564734 277538
rect 564114 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 564734 277454
rect 564114 241774 564734 277218
rect 564114 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 564734 241774
rect 564114 241454 564734 241538
rect 564114 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 564734 241454
rect 564114 205774 564734 241218
rect 564114 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 564734 205774
rect 564114 205454 564734 205538
rect 564114 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 564734 205454
rect 564114 169774 564734 205218
rect 564114 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 564734 169774
rect 564114 169454 564734 169538
rect 564114 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 564734 169454
rect 564114 133774 564734 169218
rect 564114 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 564734 133774
rect 564114 133454 564734 133538
rect 564114 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 564734 133454
rect 564114 97774 564734 133218
rect 564114 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 564734 97774
rect 564114 97454 564734 97538
rect 564114 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 564734 97454
rect 564114 61774 564734 97218
rect 564114 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 564734 61774
rect 564114 61454 564734 61538
rect 564114 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 564734 61454
rect 564114 25774 564734 61218
rect 564114 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 564734 25774
rect 564114 25454 564734 25538
rect 564114 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 564734 25454
rect 564114 -6106 564734 25218
rect 564114 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 564734 -6106
rect 564114 -6426 564734 -6342
rect 564114 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 564734 -6426
rect 564114 -7654 564734 -6662
rect 567834 711558 568454 711590
rect 567834 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 568454 711558
rect 567834 711238 568454 711322
rect 567834 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 568454 711238
rect 567834 677494 568454 711002
rect 567834 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 568454 677494
rect 567834 677174 568454 677258
rect 567834 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 568454 677174
rect 567834 641494 568454 676938
rect 567834 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 568454 641494
rect 567834 641174 568454 641258
rect 567834 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 568454 641174
rect 567834 605494 568454 640938
rect 567834 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 568454 605494
rect 567834 605174 568454 605258
rect 567834 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 568454 605174
rect 567834 569494 568454 604938
rect 567834 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 568454 569494
rect 567834 569174 568454 569258
rect 567834 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 568454 569174
rect 567834 533494 568454 568938
rect 567834 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 568454 533494
rect 567834 533174 568454 533258
rect 567834 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 568454 533174
rect 567834 497494 568454 532938
rect 567834 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 568454 497494
rect 567834 497174 568454 497258
rect 567834 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 568454 497174
rect 567834 461494 568454 496938
rect 567834 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 568454 461494
rect 567834 461174 568454 461258
rect 567834 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 568454 461174
rect 567834 425494 568454 460938
rect 567834 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 568454 425494
rect 567834 425174 568454 425258
rect 567834 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 568454 425174
rect 567834 389494 568454 424938
rect 567834 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 568454 389494
rect 567834 389174 568454 389258
rect 567834 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 568454 389174
rect 567834 353494 568454 388938
rect 567834 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 568454 353494
rect 567834 353174 568454 353258
rect 567834 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 568454 353174
rect 567834 317494 568454 352938
rect 567834 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 568454 317494
rect 567834 317174 568454 317258
rect 567834 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 568454 317174
rect 567834 281494 568454 316938
rect 567834 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 568454 281494
rect 567834 281174 568454 281258
rect 567834 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 568454 281174
rect 567834 245494 568454 280938
rect 567834 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 568454 245494
rect 567834 245174 568454 245258
rect 567834 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 568454 245174
rect 567834 209494 568454 244938
rect 567834 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 568454 209494
rect 567834 209174 568454 209258
rect 567834 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 568454 209174
rect 567834 173494 568454 208938
rect 567834 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 568454 173494
rect 567834 173174 568454 173258
rect 567834 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 568454 173174
rect 567834 137494 568454 172938
rect 567834 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 568454 137494
rect 567834 137174 568454 137258
rect 567834 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 568454 137174
rect 567834 101494 568454 136938
rect 567834 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 568454 101494
rect 567834 101174 568454 101258
rect 567834 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 568454 101174
rect 567834 65494 568454 100938
rect 567834 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 568454 65494
rect 567834 65174 568454 65258
rect 567834 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 568454 65174
rect 567834 29494 568454 64938
rect 567834 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 568454 29494
rect 567834 29174 568454 29258
rect 567834 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 568454 29174
rect 567834 -7066 568454 28938
rect 567834 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 568454 -7066
rect 567834 -7386 568454 -7302
rect 567834 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 568454 -7386
rect 567834 -7654 568454 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect 586270 690854 586890 690938
rect 586270 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect 586270 655174 586890 690618
rect 586270 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect 586270 654854 586890 654938
rect 586270 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect 586270 619174 586890 654618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 583174 586890 618618
rect 586270 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect 586270 582854 586890 582938
rect 586270 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect 586270 547174 586890 582618
rect 586270 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect 586270 546854 586890 546938
rect 586270 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect 586270 511174 586890 546618
rect 586270 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 586270 510854 586890 510938
rect 586270 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 586270 475174 586890 510618
rect 586270 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 586270 474854 586890 474938
rect 586270 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 586270 439174 586890 474618
rect 586270 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 586270 438854 586890 438938
rect 586270 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 586270 403174 586890 438618
rect 586270 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 586270 402854 586890 402938
rect 586270 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 586270 367174 586890 402618
rect 586270 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 586270 366854 586890 366938
rect 586270 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 586270 331174 586890 366618
rect 586270 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect 586270 330854 586890 330938
rect 586270 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect 586270 295174 586890 330618
rect 586270 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect 586270 294854 586890 294938
rect 586270 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect 586270 259174 586890 294618
rect 586270 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect 586270 258854 586890 258938
rect 586270 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect 586270 223174 586890 258618
rect 586270 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect 586270 222854 586890 222938
rect 586270 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect 586270 187174 586890 222618
rect 586270 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect 586270 186854 586890 186938
rect 586270 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect 586270 151174 586890 186618
rect 586270 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect 586270 150854 586890 150938
rect 586270 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect 586270 115174 586890 150618
rect 586270 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect 586270 114854 586890 114938
rect 586270 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect 586270 79174 586890 114618
rect 586270 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect 586270 78854 586890 78938
rect 586270 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect 586270 43174 586890 78618
rect 586270 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect 586270 42854 586890 42938
rect 586270 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect 586270 7174 586890 42618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 694894 587850 706202
rect 587230 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 587850 694894
rect 587230 694574 587850 694658
rect 587230 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 587850 694574
rect 587230 658894 587850 694338
rect 587230 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 587850 658894
rect 587230 658574 587850 658658
rect 587230 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 587850 658574
rect 587230 622894 587850 658338
rect 587230 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 587850 622894
rect 587230 622574 587850 622658
rect 587230 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 587850 622574
rect 587230 586894 587850 622338
rect 587230 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 587850 586894
rect 587230 586574 587850 586658
rect 587230 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 587850 586574
rect 587230 550894 587850 586338
rect 587230 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 587850 550894
rect 587230 550574 587850 550658
rect 587230 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 587850 550574
rect 587230 514894 587850 550338
rect 587230 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 587850 514894
rect 587230 514574 587850 514658
rect 587230 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 587850 514574
rect 587230 478894 587850 514338
rect 587230 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 587850 478894
rect 587230 478574 587850 478658
rect 587230 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 587850 478574
rect 587230 442894 587850 478338
rect 587230 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 587850 442894
rect 587230 442574 587850 442658
rect 587230 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 587850 442574
rect 587230 406894 587850 442338
rect 587230 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 587850 406894
rect 587230 406574 587850 406658
rect 587230 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 587850 406574
rect 587230 370894 587850 406338
rect 587230 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 587850 370894
rect 587230 370574 587850 370658
rect 587230 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 587850 370574
rect 587230 334894 587850 370338
rect 587230 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 587850 334894
rect 587230 334574 587850 334658
rect 587230 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 587850 334574
rect 587230 298894 587850 334338
rect 587230 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 587850 298894
rect 587230 298574 587850 298658
rect 587230 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 587850 298574
rect 587230 262894 587850 298338
rect 587230 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 587850 262894
rect 587230 262574 587850 262658
rect 587230 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 587850 262574
rect 587230 226894 587850 262338
rect 587230 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 587850 226894
rect 587230 226574 587850 226658
rect 587230 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 587850 226574
rect 587230 190894 587850 226338
rect 587230 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 587850 190894
rect 587230 190574 587850 190658
rect 587230 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 587850 190574
rect 587230 154894 587850 190338
rect 587230 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 587850 154894
rect 587230 154574 587850 154658
rect 587230 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 587850 154574
rect 587230 118894 587850 154338
rect 587230 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 587850 118894
rect 587230 118574 587850 118658
rect 587230 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 587850 118574
rect 587230 82894 587850 118338
rect 587230 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 587850 82894
rect 587230 82574 587850 82658
rect 587230 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 587850 82574
rect 587230 46894 587850 82338
rect 587230 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 587850 46894
rect 587230 46574 587850 46658
rect 587230 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 587850 46574
rect 587230 10894 587850 46338
rect 587230 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 587850 10894
rect 587230 10574 587850 10658
rect 587230 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 587850 10574
rect 587230 -2266 587850 10338
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 698614 588810 707162
rect 588190 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 588810 698614
rect 588190 698294 588810 698378
rect 588190 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 588810 698294
rect 588190 662614 588810 698058
rect 588190 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 588810 662614
rect 588190 662294 588810 662378
rect 588190 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 588810 662294
rect 588190 626614 588810 662058
rect 588190 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 588810 626614
rect 588190 626294 588810 626378
rect 588190 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 588810 626294
rect 588190 590614 588810 626058
rect 588190 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 588810 590614
rect 588190 590294 588810 590378
rect 588190 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 588810 590294
rect 588190 554614 588810 590058
rect 588190 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 588810 554614
rect 588190 554294 588810 554378
rect 588190 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 588810 554294
rect 588190 518614 588810 554058
rect 588190 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 588810 518614
rect 588190 518294 588810 518378
rect 588190 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 588810 518294
rect 588190 482614 588810 518058
rect 588190 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 588810 482614
rect 588190 482294 588810 482378
rect 588190 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 588810 482294
rect 588190 446614 588810 482058
rect 588190 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 588810 446614
rect 588190 446294 588810 446378
rect 588190 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 588810 446294
rect 588190 410614 588810 446058
rect 588190 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 588810 410614
rect 588190 410294 588810 410378
rect 588190 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 588810 410294
rect 588190 374614 588810 410058
rect 588190 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 588810 374614
rect 588190 374294 588810 374378
rect 588190 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 588810 374294
rect 588190 338614 588810 374058
rect 588190 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 588810 338614
rect 588190 338294 588810 338378
rect 588190 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 588810 338294
rect 588190 302614 588810 338058
rect 588190 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 588810 302614
rect 588190 302294 588810 302378
rect 588190 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 588810 302294
rect 588190 266614 588810 302058
rect 588190 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 588810 266614
rect 588190 266294 588810 266378
rect 588190 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 588810 266294
rect 588190 230614 588810 266058
rect 588190 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 588810 230614
rect 588190 230294 588810 230378
rect 588190 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 588810 230294
rect 588190 194614 588810 230058
rect 588190 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 588810 194614
rect 588190 194294 588810 194378
rect 588190 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 588810 194294
rect 588190 158614 588810 194058
rect 588190 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 588810 158614
rect 588190 158294 588810 158378
rect 588190 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 588810 158294
rect 588190 122614 588810 158058
rect 588190 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 588810 122614
rect 588190 122294 588810 122378
rect 588190 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 588810 122294
rect 588190 86614 588810 122058
rect 588190 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 588810 86614
rect 588190 86294 588810 86378
rect 588190 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 588810 86294
rect 588190 50614 588810 86058
rect 588190 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 588810 50614
rect 588190 50294 588810 50378
rect 588190 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 588810 50294
rect 588190 14614 588810 50058
rect 588190 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 588810 14614
rect 588190 14294 588810 14378
rect 588190 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 588810 14294
rect 588190 -3226 588810 14058
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 666334 589770 708122
rect 589150 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 589770 666334
rect 589150 666014 589770 666098
rect 589150 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 589770 666014
rect 589150 630334 589770 665778
rect 589150 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 589770 630334
rect 589150 630014 589770 630098
rect 589150 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 589770 630014
rect 589150 594334 589770 629778
rect 589150 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 589770 594334
rect 589150 594014 589770 594098
rect 589150 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 589770 594014
rect 589150 558334 589770 593778
rect 589150 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 589770 558334
rect 589150 558014 589770 558098
rect 589150 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 589770 558014
rect 589150 522334 589770 557778
rect 589150 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 589770 522334
rect 589150 522014 589770 522098
rect 589150 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 589770 522014
rect 589150 486334 589770 521778
rect 589150 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 589770 486334
rect 589150 486014 589770 486098
rect 589150 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 589770 486014
rect 589150 450334 589770 485778
rect 589150 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 589770 450334
rect 589150 450014 589770 450098
rect 589150 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 589770 450014
rect 589150 414334 589770 449778
rect 589150 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 589770 414334
rect 589150 414014 589770 414098
rect 589150 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 589770 414014
rect 589150 378334 589770 413778
rect 589150 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 589770 378334
rect 589150 378014 589770 378098
rect 589150 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 589770 378014
rect 589150 342334 589770 377778
rect 589150 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 589770 342334
rect 589150 342014 589770 342098
rect 589150 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 589770 342014
rect 589150 306334 589770 341778
rect 589150 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 589770 306334
rect 589150 306014 589770 306098
rect 589150 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 589770 306014
rect 589150 270334 589770 305778
rect 589150 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 589770 270334
rect 589150 270014 589770 270098
rect 589150 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 589770 270014
rect 589150 234334 589770 269778
rect 589150 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 589770 234334
rect 589150 234014 589770 234098
rect 589150 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 589770 234014
rect 589150 198334 589770 233778
rect 589150 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 589770 198334
rect 589150 198014 589770 198098
rect 589150 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 589770 198014
rect 589150 162334 589770 197778
rect 589150 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 589770 162334
rect 589150 162014 589770 162098
rect 589150 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 589770 162014
rect 589150 126334 589770 161778
rect 589150 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 589770 126334
rect 589150 126014 589770 126098
rect 589150 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 589770 126014
rect 589150 90334 589770 125778
rect 589150 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 589770 90334
rect 589150 90014 589770 90098
rect 589150 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 589770 90014
rect 589150 54334 589770 89778
rect 589150 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 589770 54334
rect 589150 54014 589770 54098
rect 589150 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 589770 54014
rect 589150 18334 589770 53778
rect 589150 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 589770 18334
rect 589150 18014 589770 18098
rect 589150 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 589770 18014
rect 589150 -4186 589770 17778
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 670054 590730 709082
rect 590110 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 590730 670054
rect 590110 669734 590730 669818
rect 590110 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 590730 669734
rect 590110 634054 590730 669498
rect 590110 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 590730 634054
rect 590110 633734 590730 633818
rect 590110 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 590730 633734
rect 590110 598054 590730 633498
rect 590110 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 590730 598054
rect 590110 597734 590730 597818
rect 590110 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 590730 597734
rect 590110 562054 590730 597498
rect 590110 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 590730 562054
rect 590110 561734 590730 561818
rect 590110 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 590730 561734
rect 590110 526054 590730 561498
rect 590110 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 590730 526054
rect 590110 525734 590730 525818
rect 590110 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 590730 525734
rect 590110 490054 590730 525498
rect 590110 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 590730 490054
rect 590110 489734 590730 489818
rect 590110 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 590730 489734
rect 590110 454054 590730 489498
rect 590110 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 590730 454054
rect 590110 453734 590730 453818
rect 590110 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 590730 453734
rect 590110 418054 590730 453498
rect 590110 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 590730 418054
rect 590110 417734 590730 417818
rect 590110 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 590730 417734
rect 590110 382054 590730 417498
rect 590110 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 590730 382054
rect 590110 381734 590730 381818
rect 590110 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 590730 381734
rect 590110 346054 590730 381498
rect 590110 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 590730 346054
rect 590110 345734 590730 345818
rect 590110 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 590730 345734
rect 590110 310054 590730 345498
rect 590110 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 590730 310054
rect 590110 309734 590730 309818
rect 590110 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 590730 309734
rect 590110 274054 590730 309498
rect 590110 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 590730 274054
rect 590110 273734 590730 273818
rect 590110 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 590730 273734
rect 590110 238054 590730 273498
rect 590110 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 590730 238054
rect 590110 237734 590730 237818
rect 590110 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 590730 237734
rect 590110 202054 590730 237498
rect 590110 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 590730 202054
rect 590110 201734 590730 201818
rect 590110 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 590730 201734
rect 590110 166054 590730 201498
rect 590110 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 590730 166054
rect 590110 165734 590730 165818
rect 590110 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 590730 165734
rect 590110 130054 590730 165498
rect 590110 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 590730 130054
rect 590110 129734 590730 129818
rect 590110 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 590730 129734
rect 590110 94054 590730 129498
rect 590110 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 590730 94054
rect 590110 93734 590730 93818
rect 590110 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 590730 93734
rect 590110 58054 590730 93498
rect 590110 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 590730 58054
rect 590110 57734 590730 57818
rect 590110 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 590730 57734
rect 590110 22054 590730 57498
rect 590110 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 590730 22054
rect 590110 21734 590730 21818
rect 590110 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 590730 21734
rect 590110 -5146 590730 21498
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 673774 591690 710042
rect 591070 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 591690 673774
rect 591070 673454 591690 673538
rect 591070 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 591690 673454
rect 591070 637774 591690 673218
rect 591070 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 591690 637774
rect 591070 637454 591690 637538
rect 591070 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 591690 637454
rect 591070 601774 591690 637218
rect 591070 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 591690 601774
rect 591070 601454 591690 601538
rect 591070 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 591690 601454
rect 591070 565774 591690 601218
rect 591070 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 591690 565774
rect 591070 565454 591690 565538
rect 591070 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 591690 565454
rect 591070 529774 591690 565218
rect 591070 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 591690 529774
rect 591070 529454 591690 529538
rect 591070 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 591690 529454
rect 591070 493774 591690 529218
rect 591070 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 591690 493774
rect 591070 493454 591690 493538
rect 591070 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 591690 493454
rect 591070 457774 591690 493218
rect 591070 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 591690 457774
rect 591070 457454 591690 457538
rect 591070 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 591690 457454
rect 591070 421774 591690 457218
rect 591070 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 591690 421774
rect 591070 421454 591690 421538
rect 591070 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 591690 421454
rect 591070 385774 591690 421218
rect 591070 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 591690 385774
rect 591070 385454 591690 385538
rect 591070 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 591690 385454
rect 591070 349774 591690 385218
rect 591070 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 591690 349774
rect 591070 349454 591690 349538
rect 591070 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 591690 349454
rect 591070 313774 591690 349218
rect 591070 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 591690 313774
rect 591070 313454 591690 313538
rect 591070 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 591690 313454
rect 591070 277774 591690 313218
rect 591070 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 591690 277774
rect 591070 277454 591690 277538
rect 591070 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 591690 277454
rect 591070 241774 591690 277218
rect 591070 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 591690 241774
rect 591070 241454 591690 241538
rect 591070 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 591690 241454
rect 591070 205774 591690 241218
rect 591070 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 591690 205774
rect 591070 205454 591690 205538
rect 591070 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 591690 205454
rect 591070 169774 591690 205218
rect 591070 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 591690 169774
rect 591070 169454 591690 169538
rect 591070 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 591690 169454
rect 591070 133774 591690 169218
rect 591070 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 591690 133774
rect 591070 133454 591690 133538
rect 591070 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 591690 133454
rect 591070 97774 591690 133218
rect 591070 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 591690 97774
rect 591070 97454 591690 97538
rect 591070 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 591690 97454
rect 591070 61774 591690 97218
rect 591070 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 591690 61774
rect 591070 61454 591690 61538
rect 591070 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 591690 61454
rect 591070 25774 591690 61218
rect 591070 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 591690 25774
rect 591070 25454 591690 25538
rect 591070 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 591690 25454
rect 591070 -6106 591690 25218
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 677494 592650 711002
rect 592030 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect 592030 677174 592650 677258
rect 592030 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect 592030 641494 592650 676938
rect 592030 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect 592030 641174 592650 641258
rect 592030 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect 592030 605494 592650 640938
rect 592030 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect 592030 605174 592650 605258
rect 592030 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect 592030 569494 592650 604938
rect 592030 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect 592030 569174 592650 569258
rect 592030 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect 592030 533494 592650 568938
rect 592030 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect 592030 533174 592650 533258
rect 592030 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect 592030 497494 592650 532938
rect 592030 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect 592030 497174 592650 497258
rect 592030 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect 592030 461494 592650 496938
rect 592030 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect 592030 461174 592650 461258
rect 592030 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect 592030 425494 592650 460938
rect 592030 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect 592030 425174 592650 425258
rect 592030 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect 592030 389494 592650 424938
rect 592030 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect 592030 389174 592650 389258
rect 592030 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect 592030 353494 592650 388938
rect 592030 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect 592030 353174 592650 353258
rect 592030 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect 592030 317494 592650 352938
rect 592030 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect 592030 317174 592650 317258
rect 592030 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect 592030 281494 592650 316938
rect 592030 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect 592030 281174 592650 281258
rect 592030 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect 592030 245494 592650 280938
rect 592030 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect 592030 245174 592650 245258
rect 592030 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect 592030 209494 592650 244938
rect 592030 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect 592030 209174 592650 209258
rect 592030 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect 592030 173494 592650 208938
rect 592030 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect 592030 173174 592650 173258
rect 592030 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect 592030 137494 592650 172938
rect 592030 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect 592030 137174 592650 137258
rect 592030 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect 592030 101494 592650 136938
rect 592030 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect 592030 101174 592650 101258
rect 592030 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect 592030 65494 592650 100938
rect 592030 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect 592030 65174 592650 65258
rect 592030 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect 592030 29494 592650 64938
rect 592030 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect 592030 29174 592650 29258
rect 592030 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect 592030 -7066 592650 28938
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 677258 -8458 677494
rect -8374 677258 -8138 677494
rect -8694 676938 -8458 677174
rect -8374 676938 -8138 677174
rect -8694 641258 -8458 641494
rect -8374 641258 -8138 641494
rect -8694 640938 -8458 641174
rect -8374 640938 -8138 641174
rect -8694 605258 -8458 605494
rect -8374 605258 -8138 605494
rect -8694 604938 -8458 605174
rect -8374 604938 -8138 605174
rect -8694 569258 -8458 569494
rect -8374 569258 -8138 569494
rect -8694 568938 -8458 569174
rect -8374 568938 -8138 569174
rect -8694 533258 -8458 533494
rect -8374 533258 -8138 533494
rect -8694 532938 -8458 533174
rect -8374 532938 -8138 533174
rect -8694 497258 -8458 497494
rect -8374 497258 -8138 497494
rect -8694 496938 -8458 497174
rect -8374 496938 -8138 497174
rect -8694 461258 -8458 461494
rect -8374 461258 -8138 461494
rect -8694 460938 -8458 461174
rect -8374 460938 -8138 461174
rect -8694 425258 -8458 425494
rect -8374 425258 -8138 425494
rect -8694 424938 -8458 425174
rect -8374 424938 -8138 425174
rect -8694 389258 -8458 389494
rect -8374 389258 -8138 389494
rect -8694 388938 -8458 389174
rect -8374 388938 -8138 389174
rect -8694 353258 -8458 353494
rect -8374 353258 -8138 353494
rect -8694 352938 -8458 353174
rect -8374 352938 -8138 353174
rect -8694 317258 -8458 317494
rect -8374 317258 -8138 317494
rect -8694 316938 -8458 317174
rect -8374 316938 -8138 317174
rect -8694 281258 -8458 281494
rect -8374 281258 -8138 281494
rect -8694 280938 -8458 281174
rect -8374 280938 -8138 281174
rect -8694 245258 -8458 245494
rect -8374 245258 -8138 245494
rect -8694 244938 -8458 245174
rect -8374 244938 -8138 245174
rect -8694 209258 -8458 209494
rect -8374 209258 -8138 209494
rect -8694 208938 -8458 209174
rect -8374 208938 -8138 209174
rect -8694 173258 -8458 173494
rect -8374 173258 -8138 173494
rect -8694 172938 -8458 173174
rect -8374 172938 -8138 173174
rect -8694 137258 -8458 137494
rect -8374 137258 -8138 137494
rect -8694 136938 -8458 137174
rect -8374 136938 -8138 137174
rect -8694 101258 -8458 101494
rect -8374 101258 -8138 101494
rect -8694 100938 -8458 101174
rect -8374 100938 -8138 101174
rect -8694 65258 -8458 65494
rect -8374 65258 -8138 65494
rect -8694 64938 -8458 65174
rect -8374 64938 -8138 65174
rect -8694 29258 -8458 29494
rect -8374 29258 -8138 29494
rect -8694 28938 -8458 29174
rect -8374 28938 -8138 29174
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 673538 -7498 673774
rect -7414 673538 -7178 673774
rect -7734 673218 -7498 673454
rect -7414 673218 -7178 673454
rect -7734 637538 -7498 637774
rect -7414 637538 -7178 637774
rect -7734 637218 -7498 637454
rect -7414 637218 -7178 637454
rect -7734 601538 -7498 601774
rect -7414 601538 -7178 601774
rect -7734 601218 -7498 601454
rect -7414 601218 -7178 601454
rect -7734 565538 -7498 565774
rect -7414 565538 -7178 565774
rect -7734 565218 -7498 565454
rect -7414 565218 -7178 565454
rect -7734 529538 -7498 529774
rect -7414 529538 -7178 529774
rect -7734 529218 -7498 529454
rect -7414 529218 -7178 529454
rect -7734 493538 -7498 493774
rect -7414 493538 -7178 493774
rect -7734 493218 -7498 493454
rect -7414 493218 -7178 493454
rect -7734 457538 -7498 457774
rect -7414 457538 -7178 457774
rect -7734 457218 -7498 457454
rect -7414 457218 -7178 457454
rect -7734 421538 -7498 421774
rect -7414 421538 -7178 421774
rect -7734 421218 -7498 421454
rect -7414 421218 -7178 421454
rect -7734 385538 -7498 385774
rect -7414 385538 -7178 385774
rect -7734 385218 -7498 385454
rect -7414 385218 -7178 385454
rect -7734 349538 -7498 349774
rect -7414 349538 -7178 349774
rect -7734 349218 -7498 349454
rect -7414 349218 -7178 349454
rect -7734 313538 -7498 313774
rect -7414 313538 -7178 313774
rect -7734 313218 -7498 313454
rect -7414 313218 -7178 313454
rect -7734 277538 -7498 277774
rect -7414 277538 -7178 277774
rect -7734 277218 -7498 277454
rect -7414 277218 -7178 277454
rect -7734 241538 -7498 241774
rect -7414 241538 -7178 241774
rect -7734 241218 -7498 241454
rect -7414 241218 -7178 241454
rect -7734 205538 -7498 205774
rect -7414 205538 -7178 205774
rect -7734 205218 -7498 205454
rect -7414 205218 -7178 205454
rect -7734 169538 -7498 169774
rect -7414 169538 -7178 169774
rect -7734 169218 -7498 169454
rect -7414 169218 -7178 169454
rect -7734 133538 -7498 133774
rect -7414 133538 -7178 133774
rect -7734 133218 -7498 133454
rect -7414 133218 -7178 133454
rect -7734 97538 -7498 97774
rect -7414 97538 -7178 97774
rect -7734 97218 -7498 97454
rect -7414 97218 -7178 97454
rect -7734 61538 -7498 61774
rect -7414 61538 -7178 61774
rect -7734 61218 -7498 61454
rect -7414 61218 -7178 61454
rect -7734 25538 -7498 25774
rect -7414 25538 -7178 25774
rect -7734 25218 -7498 25454
rect -7414 25218 -7178 25454
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 669818 -6538 670054
rect -6454 669818 -6218 670054
rect -6774 669498 -6538 669734
rect -6454 669498 -6218 669734
rect -6774 633818 -6538 634054
rect -6454 633818 -6218 634054
rect -6774 633498 -6538 633734
rect -6454 633498 -6218 633734
rect -6774 597818 -6538 598054
rect -6454 597818 -6218 598054
rect -6774 597498 -6538 597734
rect -6454 597498 -6218 597734
rect -6774 561818 -6538 562054
rect -6454 561818 -6218 562054
rect -6774 561498 -6538 561734
rect -6454 561498 -6218 561734
rect -6774 525818 -6538 526054
rect -6454 525818 -6218 526054
rect -6774 525498 -6538 525734
rect -6454 525498 -6218 525734
rect -6774 489818 -6538 490054
rect -6454 489818 -6218 490054
rect -6774 489498 -6538 489734
rect -6454 489498 -6218 489734
rect -6774 453818 -6538 454054
rect -6454 453818 -6218 454054
rect -6774 453498 -6538 453734
rect -6454 453498 -6218 453734
rect -6774 417818 -6538 418054
rect -6454 417818 -6218 418054
rect -6774 417498 -6538 417734
rect -6454 417498 -6218 417734
rect -6774 381818 -6538 382054
rect -6454 381818 -6218 382054
rect -6774 381498 -6538 381734
rect -6454 381498 -6218 381734
rect -6774 345818 -6538 346054
rect -6454 345818 -6218 346054
rect -6774 345498 -6538 345734
rect -6454 345498 -6218 345734
rect -6774 309818 -6538 310054
rect -6454 309818 -6218 310054
rect -6774 309498 -6538 309734
rect -6454 309498 -6218 309734
rect -6774 273818 -6538 274054
rect -6454 273818 -6218 274054
rect -6774 273498 -6538 273734
rect -6454 273498 -6218 273734
rect -6774 237818 -6538 238054
rect -6454 237818 -6218 238054
rect -6774 237498 -6538 237734
rect -6454 237498 -6218 237734
rect -6774 201818 -6538 202054
rect -6454 201818 -6218 202054
rect -6774 201498 -6538 201734
rect -6454 201498 -6218 201734
rect -6774 165818 -6538 166054
rect -6454 165818 -6218 166054
rect -6774 165498 -6538 165734
rect -6454 165498 -6218 165734
rect -6774 129818 -6538 130054
rect -6454 129818 -6218 130054
rect -6774 129498 -6538 129734
rect -6454 129498 -6218 129734
rect -6774 93818 -6538 94054
rect -6454 93818 -6218 94054
rect -6774 93498 -6538 93734
rect -6454 93498 -6218 93734
rect -6774 57818 -6538 58054
rect -6454 57818 -6218 58054
rect -6774 57498 -6538 57734
rect -6454 57498 -6218 57734
rect -6774 21818 -6538 22054
rect -6454 21818 -6218 22054
rect -6774 21498 -6538 21734
rect -6454 21498 -6218 21734
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 666098 -5578 666334
rect -5494 666098 -5258 666334
rect -5814 665778 -5578 666014
rect -5494 665778 -5258 666014
rect -5814 630098 -5578 630334
rect -5494 630098 -5258 630334
rect -5814 629778 -5578 630014
rect -5494 629778 -5258 630014
rect -5814 594098 -5578 594334
rect -5494 594098 -5258 594334
rect -5814 593778 -5578 594014
rect -5494 593778 -5258 594014
rect -5814 558098 -5578 558334
rect -5494 558098 -5258 558334
rect -5814 557778 -5578 558014
rect -5494 557778 -5258 558014
rect -5814 522098 -5578 522334
rect -5494 522098 -5258 522334
rect -5814 521778 -5578 522014
rect -5494 521778 -5258 522014
rect -5814 486098 -5578 486334
rect -5494 486098 -5258 486334
rect -5814 485778 -5578 486014
rect -5494 485778 -5258 486014
rect -5814 450098 -5578 450334
rect -5494 450098 -5258 450334
rect -5814 449778 -5578 450014
rect -5494 449778 -5258 450014
rect -5814 414098 -5578 414334
rect -5494 414098 -5258 414334
rect -5814 413778 -5578 414014
rect -5494 413778 -5258 414014
rect -5814 378098 -5578 378334
rect -5494 378098 -5258 378334
rect -5814 377778 -5578 378014
rect -5494 377778 -5258 378014
rect -5814 342098 -5578 342334
rect -5494 342098 -5258 342334
rect -5814 341778 -5578 342014
rect -5494 341778 -5258 342014
rect -5814 306098 -5578 306334
rect -5494 306098 -5258 306334
rect -5814 305778 -5578 306014
rect -5494 305778 -5258 306014
rect -5814 270098 -5578 270334
rect -5494 270098 -5258 270334
rect -5814 269778 -5578 270014
rect -5494 269778 -5258 270014
rect -5814 234098 -5578 234334
rect -5494 234098 -5258 234334
rect -5814 233778 -5578 234014
rect -5494 233778 -5258 234014
rect -5814 198098 -5578 198334
rect -5494 198098 -5258 198334
rect -5814 197778 -5578 198014
rect -5494 197778 -5258 198014
rect -5814 162098 -5578 162334
rect -5494 162098 -5258 162334
rect -5814 161778 -5578 162014
rect -5494 161778 -5258 162014
rect -5814 126098 -5578 126334
rect -5494 126098 -5258 126334
rect -5814 125778 -5578 126014
rect -5494 125778 -5258 126014
rect -5814 90098 -5578 90334
rect -5494 90098 -5258 90334
rect -5814 89778 -5578 90014
rect -5494 89778 -5258 90014
rect -5814 54098 -5578 54334
rect -5494 54098 -5258 54334
rect -5814 53778 -5578 54014
rect -5494 53778 -5258 54014
rect -5814 18098 -5578 18334
rect -5494 18098 -5258 18334
rect -5814 17778 -5578 18014
rect -5494 17778 -5258 18014
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 698378 -4618 698614
rect -4534 698378 -4298 698614
rect -4854 698058 -4618 698294
rect -4534 698058 -4298 698294
rect -4854 662378 -4618 662614
rect -4534 662378 -4298 662614
rect -4854 662058 -4618 662294
rect -4534 662058 -4298 662294
rect -4854 626378 -4618 626614
rect -4534 626378 -4298 626614
rect -4854 626058 -4618 626294
rect -4534 626058 -4298 626294
rect -4854 590378 -4618 590614
rect -4534 590378 -4298 590614
rect -4854 590058 -4618 590294
rect -4534 590058 -4298 590294
rect -4854 554378 -4618 554614
rect -4534 554378 -4298 554614
rect -4854 554058 -4618 554294
rect -4534 554058 -4298 554294
rect -4854 518378 -4618 518614
rect -4534 518378 -4298 518614
rect -4854 518058 -4618 518294
rect -4534 518058 -4298 518294
rect -4854 482378 -4618 482614
rect -4534 482378 -4298 482614
rect -4854 482058 -4618 482294
rect -4534 482058 -4298 482294
rect -4854 446378 -4618 446614
rect -4534 446378 -4298 446614
rect -4854 446058 -4618 446294
rect -4534 446058 -4298 446294
rect -4854 410378 -4618 410614
rect -4534 410378 -4298 410614
rect -4854 410058 -4618 410294
rect -4534 410058 -4298 410294
rect -4854 374378 -4618 374614
rect -4534 374378 -4298 374614
rect -4854 374058 -4618 374294
rect -4534 374058 -4298 374294
rect -4854 338378 -4618 338614
rect -4534 338378 -4298 338614
rect -4854 338058 -4618 338294
rect -4534 338058 -4298 338294
rect -4854 302378 -4618 302614
rect -4534 302378 -4298 302614
rect -4854 302058 -4618 302294
rect -4534 302058 -4298 302294
rect -4854 266378 -4618 266614
rect -4534 266378 -4298 266614
rect -4854 266058 -4618 266294
rect -4534 266058 -4298 266294
rect -4854 230378 -4618 230614
rect -4534 230378 -4298 230614
rect -4854 230058 -4618 230294
rect -4534 230058 -4298 230294
rect -4854 194378 -4618 194614
rect -4534 194378 -4298 194614
rect -4854 194058 -4618 194294
rect -4534 194058 -4298 194294
rect -4854 158378 -4618 158614
rect -4534 158378 -4298 158614
rect -4854 158058 -4618 158294
rect -4534 158058 -4298 158294
rect -4854 122378 -4618 122614
rect -4534 122378 -4298 122614
rect -4854 122058 -4618 122294
rect -4534 122058 -4298 122294
rect -4854 86378 -4618 86614
rect -4534 86378 -4298 86614
rect -4854 86058 -4618 86294
rect -4534 86058 -4298 86294
rect -4854 50378 -4618 50614
rect -4534 50378 -4298 50614
rect -4854 50058 -4618 50294
rect -4534 50058 -4298 50294
rect -4854 14378 -4618 14614
rect -4534 14378 -4298 14614
rect -4854 14058 -4618 14294
rect -4534 14058 -4298 14294
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 694658 -3658 694894
rect -3574 694658 -3338 694894
rect -3894 694338 -3658 694574
rect -3574 694338 -3338 694574
rect -3894 658658 -3658 658894
rect -3574 658658 -3338 658894
rect -3894 658338 -3658 658574
rect -3574 658338 -3338 658574
rect -3894 622658 -3658 622894
rect -3574 622658 -3338 622894
rect -3894 622338 -3658 622574
rect -3574 622338 -3338 622574
rect -3894 586658 -3658 586894
rect -3574 586658 -3338 586894
rect -3894 586338 -3658 586574
rect -3574 586338 -3338 586574
rect -3894 550658 -3658 550894
rect -3574 550658 -3338 550894
rect -3894 550338 -3658 550574
rect -3574 550338 -3338 550574
rect -3894 514658 -3658 514894
rect -3574 514658 -3338 514894
rect -3894 514338 -3658 514574
rect -3574 514338 -3338 514574
rect -3894 478658 -3658 478894
rect -3574 478658 -3338 478894
rect -3894 478338 -3658 478574
rect -3574 478338 -3338 478574
rect -3894 442658 -3658 442894
rect -3574 442658 -3338 442894
rect -3894 442338 -3658 442574
rect -3574 442338 -3338 442574
rect -3894 406658 -3658 406894
rect -3574 406658 -3338 406894
rect -3894 406338 -3658 406574
rect -3574 406338 -3338 406574
rect -3894 370658 -3658 370894
rect -3574 370658 -3338 370894
rect -3894 370338 -3658 370574
rect -3574 370338 -3338 370574
rect -3894 334658 -3658 334894
rect -3574 334658 -3338 334894
rect -3894 334338 -3658 334574
rect -3574 334338 -3338 334574
rect -3894 298658 -3658 298894
rect -3574 298658 -3338 298894
rect -3894 298338 -3658 298574
rect -3574 298338 -3338 298574
rect -3894 262658 -3658 262894
rect -3574 262658 -3338 262894
rect -3894 262338 -3658 262574
rect -3574 262338 -3338 262574
rect -3894 226658 -3658 226894
rect -3574 226658 -3338 226894
rect -3894 226338 -3658 226574
rect -3574 226338 -3338 226574
rect -3894 190658 -3658 190894
rect -3574 190658 -3338 190894
rect -3894 190338 -3658 190574
rect -3574 190338 -3338 190574
rect -3894 154658 -3658 154894
rect -3574 154658 -3338 154894
rect -3894 154338 -3658 154574
rect -3574 154338 -3338 154574
rect -3894 118658 -3658 118894
rect -3574 118658 -3338 118894
rect -3894 118338 -3658 118574
rect -3574 118338 -3338 118574
rect -3894 82658 -3658 82894
rect -3574 82658 -3338 82894
rect -3894 82338 -3658 82574
rect -3574 82338 -3338 82574
rect -3894 46658 -3658 46894
rect -3574 46658 -3338 46894
rect -3894 46338 -3658 46574
rect -3574 46338 -3338 46574
rect -3894 10658 -3658 10894
rect -3574 10658 -3338 10894
rect -3894 10338 -3658 10574
rect -3574 10338 -3338 10574
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 690938 -2698 691174
rect -2614 690938 -2378 691174
rect -2934 690618 -2698 690854
rect -2614 690618 -2378 690854
rect -2934 654938 -2698 655174
rect -2614 654938 -2378 655174
rect -2934 654618 -2698 654854
rect -2614 654618 -2378 654854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 582938 -2698 583174
rect -2614 582938 -2378 583174
rect -2934 582618 -2698 582854
rect -2614 582618 -2378 582854
rect -2934 546938 -2698 547174
rect -2614 546938 -2378 547174
rect -2934 546618 -2698 546854
rect -2614 546618 -2378 546854
rect -2934 510938 -2698 511174
rect -2614 510938 -2378 511174
rect -2934 510618 -2698 510854
rect -2614 510618 -2378 510854
rect -2934 474938 -2698 475174
rect -2614 474938 -2378 475174
rect -2934 474618 -2698 474854
rect -2614 474618 -2378 474854
rect -2934 438938 -2698 439174
rect -2614 438938 -2378 439174
rect -2934 438618 -2698 438854
rect -2614 438618 -2378 438854
rect -2934 402938 -2698 403174
rect -2614 402938 -2378 403174
rect -2934 402618 -2698 402854
rect -2614 402618 -2378 402854
rect -2934 366938 -2698 367174
rect -2614 366938 -2378 367174
rect -2934 366618 -2698 366854
rect -2614 366618 -2378 366854
rect -2934 330938 -2698 331174
rect -2614 330938 -2378 331174
rect -2934 330618 -2698 330854
rect -2614 330618 -2378 330854
rect -2934 294938 -2698 295174
rect -2614 294938 -2378 295174
rect -2934 294618 -2698 294854
rect -2614 294618 -2378 294854
rect -2934 258938 -2698 259174
rect -2614 258938 -2378 259174
rect -2934 258618 -2698 258854
rect -2614 258618 -2378 258854
rect -2934 222938 -2698 223174
rect -2614 222938 -2378 223174
rect -2934 222618 -2698 222854
rect -2614 222618 -2378 222854
rect -2934 186938 -2698 187174
rect -2614 186938 -2378 187174
rect -2934 186618 -2698 186854
rect -2614 186618 -2378 186854
rect -2934 150938 -2698 151174
rect -2614 150938 -2378 151174
rect -2934 150618 -2698 150854
rect -2614 150618 -2378 150854
rect -2934 114938 -2698 115174
rect -2614 114938 -2378 115174
rect -2934 114618 -2698 114854
rect -2614 114618 -2378 114854
rect -2934 78938 -2698 79174
rect -2614 78938 -2378 79174
rect -2934 78618 -2698 78854
rect -2614 78618 -2378 78854
rect -2934 42938 -2698 43174
rect -2614 42938 -2378 43174
rect -2934 42618 -2698 42854
rect -2614 42618 -2378 42854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 9266 706522 9502 706758
rect 9586 706522 9822 706758
rect 9266 706202 9502 706438
rect 9586 706202 9822 706438
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect 9266 -2502 9502 -2266
rect 9586 -2502 9822 -2266
rect 9266 -2822 9502 -2586
rect 9586 -2822 9822 -2586
rect 12986 707482 13222 707718
rect 13306 707482 13542 707718
rect 12986 707162 13222 707398
rect 13306 707162 13542 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect 12986 -3462 13222 -3226
rect 13306 -3462 13542 -3226
rect 12986 -3782 13222 -3546
rect 13306 -3782 13542 -3546
rect 16706 708442 16942 708678
rect 17026 708442 17262 708678
rect 16706 708122 16942 708358
rect 17026 708122 17262 708358
rect 16706 666098 16942 666334
rect 17026 666098 17262 666334
rect 16706 665778 16942 666014
rect 17026 665778 17262 666014
rect 16706 630098 16942 630334
rect 17026 630098 17262 630334
rect 16706 629778 16942 630014
rect 17026 629778 17262 630014
rect 16706 594098 16942 594334
rect 17026 594098 17262 594334
rect 16706 593778 16942 594014
rect 17026 593778 17262 594014
rect 16706 558098 16942 558334
rect 17026 558098 17262 558334
rect 16706 557778 16942 558014
rect 17026 557778 17262 558014
rect 16706 522098 16942 522334
rect 17026 522098 17262 522334
rect 16706 521778 16942 522014
rect 17026 521778 17262 522014
rect 16706 486098 16942 486334
rect 17026 486098 17262 486334
rect 16706 485778 16942 486014
rect 17026 485778 17262 486014
rect 16706 450098 16942 450334
rect 17026 450098 17262 450334
rect 16706 449778 16942 450014
rect 17026 449778 17262 450014
rect 16706 414098 16942 414334
rect 17026 414098 17262 414334
rect 16706 413778 16942 414014
rect 17026 413778 17262 414014
rect 16706 378098 16942 378334
rect 17026 378098 17262 378334
rect 16706 377778 16942 378014
rect 17026 377778 17262 378014
rect 16706 342098 16942 342334
rect 17026 342098 17262 342334
rect 16706 341778 16942 342014
rect 17026 341778 17262 342014
rect 16706 306098 16942 306334
rect 17026 306098 17262 306334
rect 16706 305778 16942 306014
rect 17026 305778 17262 306014
rect 16706 270098 16942 270334
rect 17026 270098 17262 270334
rect 16706 269778 16942 270014
rect 17026 269778 17262 270014
rect 16706 234098 16942 234334
rect 17026 234098 17262 234334
rect 16706 233778 16942 234014
rect 17026 233778 17262 234014
rect 16706 198098 16942 198334
rect 17026 198098 17262 198334
rect 16706 197778 16942 198014
rect 17026 197778 17262 198014
rect 16706 162098 16942 162334
rect 17026 162098 17262 162334
rect 16706 161778 16942 162014
rect 17026 161778 17262 162014
rect 16706 126098 16942 126334
rect 17026 126098 17262 126334
rect 16706 125778 16942 126014
rect 17026 125778 17262 126014
rect 16706 90098 16942 90334
rect 17026 90098 17262 90334
rect 16706 89778 16942 90014
rect 17026 89778 17262 90014
rect 16706 54098 16942 54334
rect 17026 54098 17262 54334
rect 16706 53778 16942 54014
rect 17026 53778 17262 54014
rect 16706 18098 16942 18334
rect 17026 18098 17262 18334
rect 16706 17778 16942 18014
rect 17026 17778 17262 18014
rect 16706 -4422 16942 -4186
rect 17026 -4422 17262 -4186
rect 16706 -4742 16942 -4506
rect 17026 -4742 17262 -4506
rect 20426 709402 20662 709638
rect 20746 709402 20982 709638
rect 20426 709082 20662 709318
rect 20746 709082 20982 709318
rect 20426 669818 20662 670054
rect 20746 669818 20982 670054
rect 20426 669498 20662 669734
rect 20746 669498 20982 669734
rect 20426 633818 20662 634054
rect 20746 633818 20982 634054
rect 20426 633498 20662 633734
rect 20746 633498 20982 633734
rect 20426 597818 20662 598054
rect 20746 597818 20982 598054
rect 20426 597498 20662 597734
rect 20746 597498 20982 597734
rect 20426 561818 20662 562054
rect 20746 561818 20982 562054
rect 20426 561498 20662 561734
rect 20746 561498 20982 561734
rect 20426 525818 20662 526054
rect 20746 525818 20982 526054
rect 20426 525498 20662 525734
rect 20746 525498 20982 525734
rect 20426 489818 20662 490054
rect 20746 489818 20982 490054
rect 20426 489498 20662 489734
rect 20746 489498 20982 489734
rect 20426 453818 20662 454054
rect 20746 453818 20982 454054
rect 20426 453498 20662 453734
rect 20746 453498 20982 453734
rect 20426 417818 20662 418054
rect 20746 417818 20982 418054
rect 20426 417498 20662 417734
rect 20746 417498 20982 417734
rect 20426 381818 20662 382054
rect 20746 381818 20982 382054
rect 20426 381498 20662 381734
rect 20746 381498 20982 381734
rect 20426 345818 20662 346054
rect 20746 345818 20982 346054
rect 20426 345498 20662 345734
rect 20746 345498 20982 345734
rect 20426 309818 20662 310054
rect 20746 309818 20982 310054
rect 20426 309498 20662 309734
rect 20746 309498 20982 309734
rect 20426 273818 20662 274054
rect 20746 273818 20982 274054
rect 20426 273498 20662 273734
rect 20746 273498 20982 273734
rect 20426 237818 20662 238054
rect 20746 237818 20982 238054
rect 20426 237498 20662 237734
rect 20746 237498 20982 237734
rect 20426 201818 20662 202054
rect 20746 201818 20982 202054
rect 20426 201498 20662 201734
rect 20746 201498 20982 201734
rect 20426 165818 20662 166054
rect 20746 165818 20982 166054
rect 20426 165498 20662 165734
rect 20746 165498 20982 165734
rect 20426 129818 20662 130054
rect 20746 129818 20982 130054
rect 20426 129498 20662 129734
rect 20746 129498 20982 129734
rect 20426 93818 20662 94054
rect 20746 93818 20982 94054
rect 20426 93498 20662 93734
rect 20746 93498 20982 93734
rect 20426 57818 20662 58054
rect 20746 57818 20982 58054
rect 20426 57498 20662 57734
rect 20746 57498 20982 57734
rect 20426 21818 20662 22054
rect 20746 21818 20982 22054
rect 20426 21498 20662 21734
rect 20746 21498 20982 21734
rect 20426 -5382 20662 -5146
rect 20746 -5382 20982 -5146
rect 20426 -5702 20662 -5466
rect 20746 -5702 20982 -5466
rect 24146 710362 24382 710598
rect 24466 710362 24702 710598
rect 24146 710042 24382 710278
rect 24466 710042 24702 710278
rect 24146 673538 24382 673774
rect 24466 673538 24702 673774
rect 24146 673218 24382 673454
rect 24466 673218 24702 673454
rect 24146 637538 24382 637774
rect 24466 637538 24702 637774
rect 24146 637218 24382 637454
rect 24466 637218 24702 637454
rect 24146 601538 24382 601774
rect 24466 601538 24702 601774
rect 24146 601218 24382 601454
rect 24466 601218 24702 601454
rect 24146 565538 24382 565774
rect 24466 565538 24702 565774
rect 24146 565218 24382 565454
rect 24466 565218 24702 565454
rect 24146 529538 24382 529774
rect 24466 529538 24702 529774
rect 24146 529218 24382 529454
rect 24466 529218 24702 529454
rect 24146 493538 24382 493774
rect 24466 493538 24702 493774
rect 24146 493218 24382 493454
rect 24466 493218 24702 493454
rect 24146 457538 24382 457774
rect 24466 457538 24702 457774
rect 24146 457218 24382 457454
rect 24466 457218 24702 457454
rect 24146 421538 24382 421774
rect 24466 421538 24702 421774
rect 24146 421218 24382 421454
rect 24466 421218 24702 421454
rect 24146 385538 24382 385774
rect 24466 385538 24702 385774
rect 24146 385218 24382 385454
rect 24466 385218 24702 385454
rect 24146 349538 24382 349774
rect 24466 349538 24702 349774
rect 24146 349218 24382 349454
rect 24466 349218 24702 349454
rect 24146 313538 24382 313774
rect 24466 313538 24702 313774
rect 24146 313218 24382 313454
rect 24466 313218 24702 313454
rect 24146 277538 24382 277774
rect 24466 277538 24702 277774
rect 24146 277218 24382 277454
rect 24466 277218 24702 277454
rect 24146 241538 24382 241774
rect 24466 241538 24702 241774
rect 24146 241218 24382 241454
rect 24466 241218 24702 241454
rect 24146 205538 24382 205774
rect 24466 205538 24702 205774
rect 24146 205218 24382 205454
rect 24466 205218 24702 205454
rect 24146 169538 24382 169774
rect 24466 169538 24702 169774
rect 24146 169218 24382 169454
rect 24466 169218 24702 169454
rect 24146 133538 24382 133774
rect 24466 133538 24702 133774
rect 24146 133218 24382 133454
rect 24466 133218 24702 133454
rect 24146 97538 24382 97774
rect 24466 97538 24702 97774
rect 24146 97218 24382 97454
rect 24466 97218 24702 97454
rect 24146 61538 24382 61774
rect 24466 61538 24702 61774
rect 24146 61218 24382 61454
rect 24466 61218 24702 61454
rect 24146 25538 24382 25774
rect 24466 25538 24702 25774
rect 24146 25218 24382 25454
rect 24466 25218 24702 25454
rect 24146 -6342 24382 -6106
rect 24466 -6342 24702 -6106
rect 24146 -6662 24382 -6426
rect 24466 -6662 24702 -6426
rect 27866 711322 28102 711558
rect 28186 711322 28422 711558
rect 27866 711002 28102 711238
rect 28186 711002 28422 711238
rect 27866 677258 28102 677494
rect 28186 677258 28422 677494
rect 27866 676938 28102 677174
rect 28186 676938 28422 677174
rect 27866 641258 28102 641494
rect 28186 641258 28422 641494
rect 27866 640938 28102 641174
rect 28186 640938 28422 641174
rect 27866 605258 28102 605494
rect 28186 605258 28422 605494
rect 27866 604938 28102 605174
rect 28186 604938 28422 605174
rect 27866 569258 28102 569494
rect 28186 569258 28422 569494
rect 27866 568938 28102 569174
rect 28186 568938 28422 569174
rect 27866 533258 28102 533494
rect 28186 533258 28422 533494
rect 27866 532938 28102 533174
rect 28186 532938 28422 533174
rect 27866 497258 28102 497494
rect 28186 497258 28422 497494
rect 27866 496938 28102 497174
rect 28186 496938 28422 497174
rect 27866 461258 28102 461494
rect 28186 461258 28422 461494
rect 27866 460938 28102 461174
rect 28186 460938 28422 461174
rect 27866 425258 28102 425494
rect 28186 425258 28422 425494
rect 27866 424938 28102 425174
rect 28186 424938 28422 425174
rect 27866 389258 28102 389494
rect 28186 389258 28422 389494
rect 27866 388938 28102 389174
rect 28186 388938 28422 389174
rect 27866 353258 28102 353494
rect 28186 353258 28422 353494
rect 27866 352938 28102 353174
rect 28186 352938 28422 353174
rect 27866 317258 28102 317494
rect 28186 317258 28422 317494
rect 27866 316938 28102 317174
rect 28186 316938 28422 317174
rect 27866 281258 28102 281494
rect 28186 281258 28422 281494
rect 27866 280938 28102 281174
rect 28186 280938 28422 281174
rect 27866 245258 28102 245494
rect 28186 245258 28422 245494
rect 27866 244938 28102 245174
rect 28186 244938 28422 245174
rect 27866 209258 28102 209494
rect 28186 209258 28422 209494
rect 27866 208938 28102 209174
rect 28186 208938 28422 209174
rect 27866 173258 28102 173494
rect 28186 173258 28422 173494
rect 27866 172938 28102 173174
rect 28186 172938 28422 173174
rect 27866 137258 28102 137494
rect 28186 137258 28422 137494
rect 27866 136938 28102 137174
rect 28186 136938 28422 137174
rect 27866 101258 28102 101494
rect 28186 101258 28422 101494
rect 27866 100938 28102 101174
rect 28186 100938 28422 101174
rect 27866 65258 28102 65494
rect 28186 65258 28422 65494
rect 27866 64938 28102 65174
rect 28186 64938 28422 65174
rect 27866 29258 28102 29494
rect 28186 29258 28422 29494
rect 27866 28938 28102 29174
rect 28186 28938 28422 29174
rect 27866 -7302 28102 -7066
rect 28186 -7302 28422 -7066
rect 27866 -7622 28102 -7386
rect 28186 -7622 28422 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 705562 41782 705798
rect 41866 705562 42102 705798
rect 41546 705242 41782 705478
rect 41866 705242 42102 705478
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -1542 41782 -1306
rect 41866 -1542 42102 -1306
rect 41546 -1862 41782 -1626
rect 41866 -1862 42102 -1626
rect 45266 706522 45502 706758
rect 45586 706522 45822 706758
rect 45266 706202 45502 706438
rect 45586 706202 45822 706438
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -2502 45502 -2266
rect 45586 -2502 45822 -2266
rect 45266 -2822 45502 -2586
rect 45586 -2822 45822 -2586
rect 48986 707482 49222 707718
rect 49306 707482 49542 707718
rect 48986 707162 49222 707398
rect 49306 707162 49542 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 48986 -3462 49222 -3226
rect 49306 -3462 49542 -3226
rect 48986 -3782 49222 -3546
rect 49306 -3782 49542 -3546
rect 52706 708442 52942 708678
rect 53026 708442 53262 708678
rect 52706 708122 52942 708358
rect 53026 708122 53262 708358
rect 52706 666098 52942 666334
rect 53026 666098 53262 666334
rect 52706 665778 52942 666014
rect 53026 665778 53262 666014
rect 52706 630098 52942 630334
rect 53026 630098 53262 630334
rect 52706 629778 52942 630014
rect 53026 629778 53262 630014
rect 52706 594098 52942 594334
rect 53026 594098 53262 594334
rect 52706 593778 52942 594014
rect 53026 593778 53262 594014
rect 52706 558098 52942 558334
rect 53026 558098 53262 558334
rect 52706 557778 52942 558014
rect 53026 557778 53262 558014
rect 52706 522098 52942 522334
rect 53026 522098 53262 522334
rect 52706 521778 52942 522014
rect 53026 521778 53262 522014
rect 52706 486098 52942 486334
rect 53026 486098 53262 486334
rect 52706 485778 52942 486014
rect 53026 485778 53262 486014
rect 52706 450098 52942 450334
rect 53026 450098 53262 450334
rect 52706 449778 52942 450014
rect 53026 449778 53262 450014
rect 52706 414098 52942 414334
rect 53026 414098 53262 414334
rect 52706 413778 52942 414014
rect 53026 413778 53262 414014
rect 52706 378098 52942 378334
rect 53026 378098 53262 378334
rect 52706 377778 52942 378014
rect 53026 377778 53262 378014
rect 52706 342098 52942 342334
rect 53026 342098 53262 342334
rect 52706 341778 52942 342014
rect 53026 341778 53262 342014
rect 52706 306098 52942 306334
rect 53026 306098 53262 306334
rect 52706 305778 52942 306014
rect 53026 305778 53262 306014
rect 52706 270098 52942 270334
rect 53026 270098 53262 270334
rect 52706 269778 52942 270014
rect 53026 269778 53262 270014
rect 52706 234098 52942 234334
rect 53026 234098 53262 234334
rect 52706 233778 52942 234014
rect 53026 233778 53262 234014
rect 52706 198098 52942 198334
rect 53026 198098 53262 198334
rect 52706 197778 52942 198014
rect 53026 197778 53262 198014
rect 52706 162098 52942 162334
rect 53026 162098 53262 162334
rect 52706 161778 52942 162014
rect 53026 161778 53262 162014
rect 52706 126098 52942 126334
rect 53026 126098 53262 126334
rect 52706 125778 52942 126014
rect 53026 125778 53262 126014
rect 52706 90098 52942 90334
rect 53026 90098 53262 90334
rect 52706 89778 52942 90014
rect 53026 89778 53262 90014
rect 52706 54098 52942 54334
rect 53026 54098 53262 54334
rect 52706 53778 52942 54014
rect 53026 53778 53262 54014
rect 52706 18098 52942 18334
rect 53026 18098 53262 18334
rect 52706 17778 52942 18014
rect 53026 17778 53262 18014
rect 52706 -4422 52942 -4186
rect 53026 -4422 53262 -4186
rect 52706 -4742 52942 -4506
rect 53026 -4742 53262 -4506
rect 56426 709402 56662 709638
rect 56746 709402 56982 709638
rect 56426 709082 56662 709318
rect 56746 709082 56982 709318
rect 56426 669818 56662 670054
rect 56746 669818 56982 670054
rect 56426 669498 56662 669734
rect 56746 669498 56982 669734
rect 56426 633818 56662 634054
rect 56746 633818 56982 634054
rect 56426 633498 56662 633734
rect 56746 633498 56982 633734
rect 56426 597818 56662 598054
rect 56746 597818 56982 598054
rect 56426 597498 56662 597734
rect 56746 597498 56982 597734
rect 56426 561818 56662 562054
rect 56746 561818 56982 562054
rect 56426 561498 56662 561734
rect 56746 561498 56982 561734
rect 56426 525818 56662 526054
rect 56746 525818 56982 526054
rect 56426 525498 56662 525734
rect 56746 525498 56982 525734
rect 56426 489818 56662 490054
rect 56746 489818 56982 490054
rect 56426 489498 56662 489734
rect 56746 489498 56982 489734
rect 56426 453818 56662 454054
rect 56746 453818 56982 454054
rect 56426 453498 56662 453734
rect 56746 453498 56982 453734
rect 56426 417818 56662 418054
rect 56746 417818 56982 418054
rect 56426 417498 56662 417734
rect 56746 417498 56982 417734
rect 56426 381818 56662 382054
rect 56746 381818 56982 382054
rect 56426 381498 56662 381734
rect 56746 381498 56982 381734
rect 56426 345818 56662 346054
rect 56746 345818 56982 346054
rect 56426 345498 56662 345734
rect 56746 345498 56982 345734
rect 56426 309818 56662 310054
rect 56746 309818 56982 310054
rect 56426 309498 56662 309734
rect 56746 309498 56982 309734
rect 56426 273818 56662 274054
rect 56746 273818 56982 274054
rect 56426 273498 56662 273734
rect 56746 273498 56982 273734
rect 56426 237818 56662 238054
rect 56746 237818 56982 238054
rect 56426 237498 56662 237734
rect 56746 237498 56982 237734
rect 56426 201818 56662 202054
rect 56746 201818 56982 202054
rect 56426 201498 56662 201734
rect 56746 201498 56982 201734
rect 56426 165818 56662 166054
rect 56746 165818 56982 166054
rect 56426 165498 56662 165734
rect 56746 165498 56982 165734
rect 56426 129818 56662 130054
rect 56746 129818 56982 130054
rect 56426 129498 56662 129734
rect 56746 129498 56982 129734
rect 56426 93818 56662 94054
rect 56746 93818 56982 94054
rect 56426 93498 56662 93734
rect 56746 93498 56982 93734
rect 56426 57818 56662 58054
rect 56746 57818 56982 58054
rect 56426 57498 56662 57734
rect 56746 57498 56982 57734
rect 56426 21818 56662 22054
rect 56746 21818 56982 22054
rect 56426 21498 56662 21734
rect 56746 21498 56982 21734
rect 56426 -5382 56662 -5146
rect 56746 -5382 56982 -5146
rect 56426 -5702 56662 -5466
rect 56746 -5702 56982 -5466
rect 60146 710362 60382 710598
rect 60466 710362 60702 710598
rect 60146 710042 60382 710278
rect 60466 710042 60702 710278
rect 60146 673538 60382 673774
rect 60466 673538 60702 673774
rect 60146 673218 60382 673454
rect 60466 673218 60702 673454
rect 60146 637538 60382 637774
rect 60466 637538 60702 637774
rect 60146 637218 60382 637454
rect 60466 637218 60702 637454
rect 60146 601538 60382 601774
rect 60466 601538 60702 601774
rect 60146 601218 60382 601454
rect 60466 601218 60702 601454
rect 60146 565538 60382 565774
rect 60466 565538 60702 565774
rect 60146 565218 60382 565454
rect 60466 565218 60702 565454
rect 60146 529538 60382 529774
rect 60466 529538 60702 529774
rect 60146 529218 60382 529454
rect 60466 529218 60702 529454
rect 60146 493538 60382 493774
rect 60466 493538 60702 493774
rect 60146 493218 60382 493454
rect 60466 493218 60702 493454
rect 60146 457538 60382 457774
rect 60466 457538 60702 457774
rect 60146 457218 60382 457454
rect 60466 457218 60702 457454
rect 60146 421538 60382 421774
rect 60466 421538 60702 421774
rect 60146 421218 60382 421454
rect 60466 421218 60702 421454
rect 60146 385538 60382 385774
rect 60466 385538 60702 385774
rect 60146 385218 60382 385454
rect 60466 385218 60702 385454
rect 60146 349538 60382 349774
rect 60466 349538 60702 349774
rect 60146 349218 60382 349454
rect 60466 349218 60702 349454
rect 60146 313538 60382 313774
rect 60466 313538 60702 313774
rect 60146 313218 60382 313454
rect 60466 313218 60702 313454
rect 60146 277538 60382 277774
rect 60466 277538 60702 277774
rect 60146 277218 60382 277454
rect 60466 277218 60702 277454
rect 60146 241538 60382 241774
rect 60466 241538 60702 241774
rect 60146 241218 60382 241454
rect 60466 241218 60702 241454
rect 60146 205538 60382 205774
rect 60466 205538 60702 205774
rect 60146 205218 60382 205454
rect 60466 205218 60702 205454
rect 60146 169538 60382 169774
rect 60466 169538 60702 169774
rect 60146 169218 60382 169454
rect 60466 169218 60702 169454
rect 60146 133538 60382 133774
rect 60466 133538 60702 133774
rect 60146 133218 60382 133454
rect 60466 133218 60702 133454
rect 60146 97538 60382 97774
rect 60466 97538 60702 97774
rect 60146 97218 60382 97454
rect 60466 97218 60702 97454
rect 60146 61538 60382 61774
rect 60466 61538 60702 61774
rect 60146 61218 60382 61454
rect 60466 61218 60702 61454
rect 60146 25538 60382 25774
rect 60466 25538 60702 25774
rect 60146 25218 60382 25454
rect 60466 25218 60702 25454
rect 60146 -6342 60382 -6106
rect 60466 -6342 60702 -6106
rect 60146 -6662 60382 -6426
rect 60466 -6662 60702 -6426
rect 63866 711322 64102 711558
rect 64186 711322 64422 711558
rect 63866 711002 64102 711238
rect 64186 711002 64422 711238
rect 63866 677258 64102 677494
rect 64186 677258 64422 677494
rect 63866 676938 64102 677174
rect 64186 676938 64422 677174
rect 63866 641258 64102 641494
rect 64186 641258 64422 641494
rect 63866 640938 64102 641174
rect 64186 640938 64422 641174
rect 63866 605258 64102 605494
rect 64186 605258 64422 605494
rect 63866 604938 64102 605174
rect 64186 604938 64422 605174
rect 63866 569258 64102 569494
rect 64186 569258 64422 569494
rect 63866 568938 64102 569174
rect 64186 568938 64422 569174
rect 63866 533258 64102 533494
rect 64186 533258 64422 533494
rect 63866 532938 64102 533174
rect 64186 532938 64422 533174
rect 63866 497258 64102 497494
rect 64186 497258 64422 497494
rect 63866 496938 64102 497174
rect 64186 496938 64422 497174
rect 63866 461258 64102 461494
rect 64186 461258 64422 461494
rect 63866 460938 64102 461174
rect 64186 460938 64422 461174
rect 63866 425258 64102 425494
rect 64186 425258 64422 425494
rect 63866 424938 64102 425174
rect 64186 424938 64422 425174
rect 63866 389258 64102 389494
rect 64186 389258 64422 389494
rect 63866 388938 64102 389174
rect 64186 388938 64422 389174
rect 63866 353258 64102 353494
rect 64186 353258 64422 353494
rect 63866 352938 64102 353174
rect 64186 352938 64422 353174
rect 63866 317258 64102 317494
rect 64186 317258 64422 317494
rect 63866 316938 64102 317174
rect 64186 316938 64422 317174
rect 63866 281258 64102 281494
rect 64186 281258 64422 281494
rect 63866 280938 64102 281174
rect 64186 280938 64422 281174
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 63866 245258 64102 245494
rect 64186 245258 64422 245494
rect 63866 244938 64102 245174
rect 64186 244938 64422 245174
rect 63866 209258 64102 209494
rect 64186 209258 64422 209494
rect 63866 208938 64102 209174
rect 64186 208938 64422 209174
rect 63866 173258 64102 173494
rect 64186 173258 64422 173494
rect 63866 172938 64102 173174
rect 64186 172938 64422 173174
rect 63866 137258 64102 137494
rect 64186 137258 64422 137494
rect 63866 136938 64102 137174
rect 64186 136938 64422 137174
rect 63866 101258 64102 101494
rect 64186 101258 64422 101494
rect 63866 100938 64102 101174
rect 64186 100938 64422 101174
rect 77546 705562 77782 705798
rect 77866 705562 78102 705798
rect 77546 705242 77782 705478
rect 77866 705242 78102 705478
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 74250 219218 74486 219454
rect 74250 218898 74486 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 81266 706522 81502 706758
rect 81586 706522 81822 706758
rect 81266 706202 81502 706438
rect 81586 706202 81822 706438
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 63866 65258 64102 65494
rect 64186 65258 64422 65494
rect 63866 64938 64102 65174
rect 64186 64938 64422 65174
rect 63866 29258 64102 29494
rect 64186 29258 64422 29494
rect 63866 28938 64102 29174
rect 64186 28938 64422 29174
rect 63866 -7302 64102 -7066
rect 64186 -7302 64422 -7066
rect 63866 -7622 64102 -7386
rect 64186 -7622 64422 -7386
rect 75206 75218 75442 75454
rect 75206 74898 75442 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 79426 78938 79662 79174
rect 79426 78618 79662 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -1542 77782 -1306
rect 77866 -1542 78102 -1306
rect 77546 -1862 77782 -1626
rect 77866 -1862 78102 -1626
rect 84986 707482 85222 707718
rect 85306 707482 85542 707718
rect 84986 707162 85222 707398
rect 85306 707162 85542 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 88706 708442 88942 708678
rect 89026 708442 89262 708678
rect 88706 708122 88942 708358
rect 89026 708122 89262 708358
rect 88706 666098 88942 666334
rect 89026 666098 89262 666334
rect 88706 665778 88942 666014
rect 89026 665778 89262 666014
rect 88706 630098 88942 630334
rect 89026 630098 89262 630334
rect 88706 629778 88942 630014
rect 89026 629778 89262 630014
rect 88706 594098 88942 594334
rect 89026 594098 89262 594334
rect 88706 593778 88942 594014
rect 89026 593778 89262 594014
rect 88706 558098 88942 558334
rect 89026 558098 89262 558334
rect 88706 557778 88942 558014
rect 89026 557778 89262 558014
rect 88706 522098 88942 522334
rect 89026 522098 89262 522334
rect 88706 521778 88942 522014
rect 89026 521778 89262 522014
rect 88706 486098 88942 486334
rect 89026 486098 89262 486334
rect 88706 485778 88942 486014
rect 89026 485778 89262 486014
rect 88706 450098 88942 450334
rect 89026 450098 89262 450334
rect 88706 449778 88942 450014
rect 89026 449778 89262 450014
rect 88706 414098 88942 414334
rect 89026 414098 89262 414334
rect 88706 413778 88942 414014
rect 89026 413778 89262 414014
rect 88706 378098 88942 378334
rect 89026 378098 89262 378334
rect 88706 377778 88942 378014
rect 89026 377778 89262 378014
rect 88706 342098 88942 342334
rect 89026 342098 89262 342334
rect 88706 341778 88942 342014
rect 89026 341778 89262 342014
rect 88706 306098 88942 306334
rect 89026 306098 89262 306334
rect 88706 305778 88942 306014
rect 89026 305778 89262 306014
rect 88706 270098 88942 270334
rect 89026 270098 89262 270334
rect 88706 269778 88942 270014
rect 89026 269778 89262 270014
rect 92426 709402 92662 709638
rect 92746 709402 92982 709638
rect 92426 709082 92662 709318
rect 92746 709082 92982 709318
rect 92426 669818 92662 670054
rect 92746 669818 92982 670054
rect 92426 669498 92662 669734
rect 92746 669498 92982 669734
rect 92426 633818 92662 634054
rect 92746 633818 92982 634054
rect 92426 633498 92662 633734
rect 92746 633498 92982 633734
rect 92426 597818 92662 598054
rect 92746 597818 92982 598054
rect 92426 597498 92662 597734
rect 92746 597498 92982 597734
rect 92426 561818 92662 562054
rect 92746 561818 92982 562054
rect 92426 561498 92662 561734
rect 92746 561498 92982 561734
rect 92426 525818 92662 526054
rect 92746 525818 92982 526054
rect 92426 525498 92662 525734
rect 92746 525498 92982 525734
rect 92426 489818 92662 490054
rect 92746 489818 92982 490054
rect 92426 489498 92662 489734
rect 92746 489498 92982 489734
rect 92426 453818 92662 454054
rect 92746 453818 92982 454054
rect 92426 453498 92662 453734
rect 92746 453498 92982 453734
rect 92426 417818 92662 418054
rect 92746 417818 92982 418054
rect 92426 417498 92662 417734
rect 92746 417498 92982 417734
rect 92426 381818 92662 382054
rect 92746 381818 92982 382054
rect 92426 381498 92662 381734
rect 92746 381498 92982 381734
rect 92426 345818 92662 346054
rect 92746 345818 92982 346054
rect 92426 345498 92662 345734
rect 92746 345498 92982 345734
rect 92426 309818 92662 310054
rect 92746 309818 92982 310054
rect 92426 309498 92662 309734
rect 92746 309498 92982 309734
rect 92426 273818 92662 274054
rect 92746 273818 92982 274054
rect 92426 273498 92662 273734
rect 92746 273498 92982 273734
rect 96146 710362 96382 710598
rect 96466 710362 96702 710598
rect 96146 710042 96382 710278
rect 96466 710042 96702 710278
rect 96146 673538 96382 673774
rect 96466 673538 96702 673774
rect 96146 673218 96382 673454
rect 96466 673218 96702 673454
rect 96146 637538 96382 637774
rect 96466 637538 96702 637774
rect 96146 637218 96382 637454
rect 96466 637218 96702 637454
rect 96146 601538 96382 601774
rect 96466 601538 96702 601774
rect 96146 601218 96382 601454
rect 96466 601218 96702 601454
rect 96146 565538 96382 565774
rect 96466 565538 96702 565774
rect 96146 565218 96382 565454
rect 96466 565218 96702 565454
rect 96146 529538 96382 529774
rect 96466 529538 96702 529774
rect 96146 529218 96382 529454
rect 96466 529218 96702 529454
rect 96146 493538 96382 493774
rect 96466 493538 96702 493774
rect 96146 493218 96382 493454
rect 96466 493218 96702 493454
rect 96146 457538 96382 457774
rect 96466 457538 96702 457774
rect 96146 457218 96382 457454
rect 96466 457218 96702 457454
rect 96146 421538 96382 421774
rect 96466 421538 96702 421774
rect 96146 421218 96382 421454
rect 96466 421218 96702 421454
rect 96146 385538 96382 385774
rect 96466 385538 96702 385774
rect 96146 385218 96382 385454
rect 96466 385218 96702 385454
rect 96146 349538 96382 349774
rect 96466 349538 96702 349774
rect 96146 349218 96382 349454
rect 96466 349218 96702 349454
rect 96146 313538 96382 313774
rect 96466 313538 96702 313774
rect 96146 313218 96382 313454
rect 96466 313218 96702 313454
rect 96146 277538 96382 277774
rect 96466 277538 96702 277774
rect 96146 277218 96382 277454
rect 96466 277218 96702 277454
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 96146 241538 96382 241774
rect 96466 241538 96702 241774
rect 96146 241218 96382 241454
rect 96466 241218 96702 241454
rect 89610 222938 89846 223174
rect 89610 222618 89846 222854
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 83647 75218 83883 75454
rect 83647 74898 83883 75134
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -2502 81502 -2266
rect 81586 -2502 81822 -2266
rect 81266 -2822 81502 -2586
rect 81586 -2822 81822 -2586
rect 88706 198098 88942 198334
rect 89026 198098 89262 198334
rect 88706 197778 88942 198014
rect 89026 197778 89262 198014
rect 88706 162098 88942 162334
rect 89026 162098 89262 162334
rect 88706 161778 88942 162014
rect 89026 161778 89262 162014
rect 88706 126098 88942 126334
rect 89026 126098 89262 126334
rect 88706 125778 88942 126014
rect 89026 125778 89262 126014
rect 92426 201818 92662 202054
rect 92746 201818 92982 202054
rect 92426 201498 92662 201734
rect 92746 201498 92982 201734
rect 92426 165818 92662 166054
rect 92746 165818 92982 166054
rect 92426 165498 92662 165734
rect 92746 165498 92982 165734
rect 92426 129818 92662 130054
rect 92746 129818 92982 130054
rect 92426 129498 92662 129734
rect 92746 129498 92982 129734
rect 96146 205538 96382 205774
rect 96466 205538 96702 205774
rect 96146 205218 96382 205454
rect 96466 205218 96702 205454
rect 96146 169538 96382 169774
rect 96466 169538 96702 169774
rect 96146 169218 96382 169454
rect 96466 169218 96702 169454
rect 96146 133538 96382 133774
rect 96466 133538 96702 133774
rect 96146 133218 96382 133454
rect 96466 133218 96702 133454
rect 99866 711322 100102 711558
rect 100186 711322 100422 711558
rect 99866 711002 100102 711238
rect 100186 711002 100422 711238
rect 99866 677258 100102 677494
rect 100186 677258 100422 677494
rect 99866 676938 100102 677174
rect 100186 676938 100422 677174
rect 99866 641258 100102 641494
rect 100186 641258 100422 641494
rect 99866 640938 100102 641174
rect 100186 640938 100422 641174
rect 99866 605258 100102 605494
rect 100186 605258 100422 605494
rect 99866 604938 100102 605174
rect 100186 604938 100422 605174
rect 99866 569258 100102 569494
rect 100186 569258 100422 569494
rect 99866 568938 100102 569174
rect 100186 568938 100422 569174
rect 99866 533258 100102 533494
rect 100186 533258 100422 533494
rect 99866 532938 100102 533174
rect 100186 532938 100422 533174
rect 99866 497258 100102 497494
rect 100186 497258 100422 497494
rect 99866 496938 100102 497174
rect 100186 496938 100422 497174
rect 99866 461258 100102 461494
rect 100186 461258 100422 461494
rect 99866 460938 100102 461174
rect 100186 460938 100422 461174
rect 99866 425258 100102 425494
rect 100186 425258 100422 425494
rect 99866 424938 100102 425174
rect 100186 424938 100422 425174
rect 99866 389258 100102 389494
rect 100186 389258 100422 389494
rect 99866 388938 100102 389174
rect 100186 388938 100422 389174
rect 99866 353258 100102 353494
rect 100186 353258 100422 353494
rect 99866 352938 100102 353174
rect 100186 352938 100422 353174
rect 99866 317258 100102 317494
rect 100186 317258 100422 317494
rect 99866 316938 100102 317174
rect 100186 316938 100422 317174
rect 99866 281258 100102 281494
rect 100186 281258 100422 281494
rect 99866 280938 100102 281174
rect 100186 280938 100422 281174
rect 99866 245258 100102 245494
rect 100186 245258 100422 245494
rect 99866 244938 100102 245174
rect 100186 244938 100422 245174
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 104970 219218 105206 219454
rect 104970 218898 105206 219134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 99866 209258 100102 209494
rect 100186 209258 100422 209494
rect 99866 208938 100102 209174
rect 100186 208938 100422 209174
rect 99866 173258 100102 173494
rect 100186 173258 100422 173494
rect 99866 172938 100102 173174
rect 100186 172938 100422 173174
rect 99866 137258 100102 137494
rect 100186 137258 100422 137494
rect 99866 136938 100102 137174
rect 100186 136938 100422 137174
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 88706 90098 88942 90334
rect 89026 90098 89262 90334
rect 88706 89778 88942 90014
rect 89026 89778 89262 90014
rect 87867 78938 88103 79174
rect 87867 78618 88103 78854
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 84986 -3462 85222 -3226
rect 85306 -3462 85542 -3226
rect 84986 -3782 85222 -3546
rect 85306 -3782 85542 -3546
rect 96308 78938 96544 79174
rect 96308 78618 96544 78854
rect 104749 78938 104985 79174
rect 104749 78618 104985 78854
rect 92088 75218 92324 75454
rect 92088 74898 92324 75134
rect 100529 75218 100765 75454
rect 100529 74898 100765 75134
rect 88706 54098 88942 54334
rect 89026 54098 89262 54334
rect 88706 53778 88942 54014
rect 89026 53778 89262 54014
rect 88706 18098 88942 18334
rect 89026 18098 89262 18334
rect 88706 17778 88942 18014
rect 89026 17778 89262 18014
rect 88706 -4422 88942 -4186
rect 89026 -4422 89262 -4186
rect 88706 -4742 88942 -4506
rect 89026 -4742 89262 -4506
rect 92426 57818 92662 58054
rect 92746 57818 92982 58054
rect 92426 57498 92662 57734
rect 92746 57498 92982 57734
rect 92426 21818 92662 22054
rect 92746 21818 92982 22054
rect 92426 21498 92662 21734
rect 92746 21498 92982 21734
rect 92426 -5382 92662 -5146
rect 92746 -5382 92982 -5146
rect 92426 -5702 92662 -5466
rect 92746 -5702 92982 -5466
rect 96146 61538 96382 61774
rect 96466 61538 96702 61774
rect 96146 61218 96382 61454
rect 96466 61218 96702 61454
rect 96146 25538 96382 25774
rect 96466 25538 96702 25774
rect 96146 25218 96382 25454
rect 96466 25218 96702 25454
rect 96146 -6342 96382 -6106
rect 96466 -6342 96702 -6106
rect 96146 -6662 96382 -6426
rect 96466 -6662 96702 -6426
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 99866 65258 100102 65494
rect 100186 65258 100422 65494
rect 99866 64938 100102 65174
rect 100186 64938 100422 65174
rect 99866 29258 100102 29494
rect 100186 29258 100422 29494
rect 99866 28938 100102 29174
rect 100186 28938 100422 29174
rect 99866 -7302 100102 -7066
rect 100186 -7302 100422 -7066
rect 99866 -7622 100102 -7386
rect 100186 -7622 100422 -7386
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 705562 113782 705798
rect 113866 705562 114102 705798
rect 113546 705242 113782 705478
rect 113866 705242 114102 705478
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -1542 113782 -1306
rect 113866 -1542 114102 -1306
rect 113546 -1862 113782 -1626
rect 113866 -1862 114102 -1626
rect 117266 706522 117502 706758
rect 117586 706522 117822 706758
rect 117266 706202 117502 706438
rect 117586 706202 117822 706438
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 120986 707482 121222 707718
rect 121306 707482 121542 707718
rect 120986 707162 121222 707398
rect 121306 707162 121542 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 124706 708442 124942 708678
rect 125026 708442 125262 708678
rect 124706 708122 124942 708358
rect 125026 708122 125262 708358
rect 124706 666098 124942 666334
rect 125026 666098 125262 666334
rect 124706 665778 124942 666014
rect 125026 665778 125262 666014
rect 124706 630098 124942 630334
rect 125026 630098 125262 630334
rect 124706 629778 124942 630014
rect 125026 629778 125262 630014
rect 124706 594098 124942 594334
rect 125026 594098 125262 594334
rect 124706 593778 124942 594014
rect 125026 593778 125262 594014
rect 124706 558098 124942 558334
rect 125026 558098 125262 558334
rect 124706 557778 124942 558014
rect 125026 557778 125262 558014
rect 124706 522098 124942 522334
rect 125026 522098 125262 522334
rect 124706 521778 124942 522014
rect 125026 521778 125262 522014
rect 124706 486098 124942 486334
rect 125026 486098 125262 486334
rect 124706 485778 124942 486014
rect 125026 485778 125262 486014
rect 124706 450098 124942 450334
rect 125026 450098 125262 450334
rect 124706 449778 124942 450014
rect 125026 449778 125262 450014
rect 124706 414098 124942 414334
rect 125026 414098 125262 414334
rect 124706 413778 124942 414014
rect 125026 413778 125262 414014
rect 124706 378098 124942 378334
rect 125026 378098 125262 378334
rect 124706 377778 124942 378014
rect 125026 377778 125262 378014
rect 124706 342098 124942 342334
rect 125026 342098 125262 342334
rect 124706 341778 124942 342014
rect 125026 341778 125262 342014
rect 124706 306098 124942 306334
rect 125026 306098 125262 306334
rect 124706 305778 124942 306014
rect 125026 305778 125262 306014
rect 124706 270098 124942 270334
rect 125026 270098 125262 270334
rect 124706 269778 124942 270014
rect 125026 269778 125262 270014
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 124706 234098 124942 234334
rect 125026 234098 125262 234334
rect 124706 233778 124942 234014
rect 125026 233778 125262 234014
rect 124706 198098 124942 198334
rect 125026 198098 125262 198334
rect 124706 197778 124942 198014
rect 125026 197778 125262 198014
rect 124706 162098 124942 162334
rect 125026 162098 125262 162334
rect 124706 161778 124942 162014
rect 125026 161778 125262 162014
rect 124706 126098 124942 126334
rect 125026 126098 125262 126334
rect 124706 125778 124942 126014
rect 125026 125778 125262 126014
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -2502 117502 -2266
rect 117586 -2502 117822 -2266
rect 117266 -2822 117502 -2586
rect 117586 -2822 117822 -2586
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 120986 -3462 121222 -3226
rect 121306 -3462 121542 -3226
rect 120986 -3782 121222 -3546
rect 121306 -3782 121542 -3546
rect 124706 90098 124942 90334
rect 125026 90098 125262 90334
rect 124706 89778 124942 90014
rect 125026 89778 125262 90014
rect 124706 54098 124942 54334
rect 125026 54098 125262 54334
rect 124706 53778 124942 54014
rect 125026 53778 125262 54014
rect 124706 18098 124942 18334
rect 125026 18098 125262 18334
rect 124706 17778 124942 18014
rect 125026 17778 125262 18014
rect 124706 -4422 124942 -4186
rect 125026 -4422 125262 -4186
rect 124706 -4742 124942 -4506
rect 125026 -4742 125262 -4506
rect 128426 709402 128662 709638
rect 128746 709402 128982 709638
rect 128426 709082 128662 709318
rect 128746 709082 128982 709318
rect 128426 669818 128662 670054
rect 128746 669818 128982 670054
rect 128426 669498 128662 669734
rect 128746 669498 128982 669734
rect 128426 633818 128662 634054
rect 128746 633818 128982 634054
rect 128426 633498 128662 633734
rect 128746 633498 128982 633734
rect 128426 597818 128662 598054
rect 128746 597818 128982 598054
rect 128426 597498 128662 597734
rect 128746 597498 128982 597734
rect 128426 561818 128662 562054
rect 128746 561818 128982 562054
rect 128426 561498 128662 561734
rect 128746 561498 128982 561734
rect 128426 525818 128662 526054
rect 128746 525818 128982 526054
rect 128426 525498 128662 525734
rect 128746 525498 128982 525734
rect 128426 489818 128662 490054
rect 128746 489818 128982 490054
rect 128426 489498 128662 489734
rect 128746 489498 128982 489734
rect 128426 453818 128662 454054
rect 128746 453818 128982 454054
rect 128426 453498 128662 453734
rect 128746 453498 128982 453734
rect 128426 417818 128662 418054
rect 128746 417818 128982 418054
rect 128426 417498 128662 417734
rect 128746 417498 128982 417734
rect 128426 381818 128662 382054
rect 128746 381818 128982 382054
rect 128426 381498 128662 381734
rect 128746 381498 128982 381734
rect 128426 345818 128662 346054
rect 128746 345818 128982 346054
rect 128426 345498 128662 345734
rect 128746 345498 128982 345734
rect 128426 309818 128662 310054
rect 128746 309818 128982 310054
rect 128426 309498 128662 309734
rect 128746 309498 128982 309734
rect 128426 273818 128662 274054
rect 128746 273818 128982 274054
rect 128426 273498 128662 273734
rect 128746 273498 128982 273734
rect 128426 237818 128662 238054
rect 128746 237818 128982 238054
rect 128426 237498 128662 237734
rect 128746 237498 128982 237734
rect 128426 201818 128662 202054
rect 128746 201818 128982 202054
rect 128426 201498 128662 201734
rect 128746 201498 128982 201734
rect 128426 165818 128662 166054
rect 128746 165818 128982 166054
rect 128426 165498 128662 165734
rect 128746 165498 128982 165734
rect 128426 129818 128662 130054
rect 128746 129818 128982 130054
rect 128426 129498 128662 129734
rect 128746 129498 128982 129734
rect 128426 93818 128662 94054
rect 128746 93818 128982 94054
rect 128426 93498 128662 93734
rect 128746 93498 128982 93734
rect 128426 57818 128662 58054
rect 128746 57818 128982 58054
rect 128426 57498 128662 57734
rect 128746 57498 128982 57734
rect 128426 21818 128662 22054
rect 128746 21818 128982 22054
rect 128426 21498 128662 21734
rect 128746 21498 128982 21734
rect 128426 -5382 128662 -5146
rect 128746 -5382 128982 -5146
rect 128426 -5702 128662 -5466
rect 128746 -5702 128982 -5466
rect 132146 710362 132382 710598
rect 132466 710362 132702 710598
rect 132146 710042 132382 710278
rect 132466 710042 132702 710278
rect 132146 673538 132382 673774
rect 132466 673538 132702 673774
rect 132146 673218 132382 673454
rect 132466 673218 132702 673454
rect 132146 637538 132382 637774
rect 132466 637538 132702 637774
rect 132146 637218 132382 637454
rect 132466 637218 132702 637454
rect 132146 601538 132382 601774
rect 132466 601538 132702 601774
rect 132146 601218 132382 601454
rect 132466 601218 132702 601454
rect 132146 565538 132382 565774
rect 132466 565538 132702 565774
rect 132146 565218 132382 565454
rect 132466 565218 132702 565454
rect 132146 529538 132382 529774
rect 132466 529538 132702 529774
rect 132146 529218 132382 529454
rect 132466 529218 132702 529454
rect 132146 493538 132382 493774
rect 132466 493538 132702 493774
rect 132146 493218 132382 493454
rect 132466 493218 132702 493454
rect 132146 457538 132382 457774
rect 132466 457538 132702 457774
rect 132146 457218 132382 457454
rect 132466 457218 132702 457454
rect 132146 421538 132382 421774
rect 132466 421538 132702 421774
rect 132146 421218 132382 421454
rect 132466 421218 132702 421454
rect 132146 385538 132382 385774
rect 132466 385538 132702 385774
rect 132146 385218 132382 385454
rect 132466 385218 132702 385454
rect 132146 349538 132382 349774
rect 132466 349538 132702 349774
rect 132146 349218 132382 349454
rect 132466 349218 132702 349454
rect 132146 313538 132382 313774
rect 132466 313538 132702 313774
rect 132146 313218 132382 313454
rect 132466 313218 132702 313454
rect 132146 277538 132382 277774
rect 132466 277538 132702 277774
rect 132146 277218 132382 277454
rect 132466 277218 132702 277454
rect 132146 241538 132382 241774
rect 132466 241538 132702 241774
rect 132146 241218 132382 241454
rect 132466 241218 132702 241454
rect 132146 205538 132382 205774
rect 132466 205538 132702 205774
rect 132146 205218 132382 205454
rect 132466 205218 132702 205454
rect 132146 169538 132382 169774
rect 132466 169538 132702 169774
rect 132146 169218 132382 169454
rect 132466 169218 132702 169454
rect 132146 133538 132382 133774
rect 132466 133538 132702 133774
rect 132146 133218 132382 133454
rect 132466 133218 132702 133454
rect 132146 97538 132382 97774
rect 132466 97538 132702 97774
rect 132146 97218 132382 97454
rect 132466 97218 132702 97454
rect 132146 61538 132382 61774
rect 132466 61538 132702 61774
rect 132146 61218 132382 61454
rect 132466 61218 132702 61454
rect 132146 25538 132382 25774
rect 132466 25538 132702 25774
rect 132146 25218 132382 25454
rect 132466 25218 132702 25454
rect 132146 -6342 132382 -6106
rect 132466 -6342 132702 -6106
rect 132146 -6662 132382 -6426
rect 132466 -6662 132702 -6426
rect 135866 711322 136102 711558
rect 136186 711322 136422 711558
rect 135866 711002 136102 711238
rect 136186 711002 136422 711238
rect 135866 677258 136102 677494
rect 136186 677258 136422 677494
rect 135866 676938 136102 677174
rect 136186 676938 136422 677174
rect 135866 641258 136102 641494
rect 136186 641258 136422 641494
rect 135866 640938 136102 641174
rect 136186 640938 136422 641174
rect 135866 605258 136102 605494
rect 136186 605258 136422 605494
rect 135866 604938 136102 605174
rect 136186 604938 136422 605174
rect 135866 569258 136102 569494
rect 136186 569258 136422 569494
rect 135866 568938 136102 569174
rect 136186 568938 136422 569174
rect 135866 533258 136102 533494
rect 136186 533258 136422 533494
rect 135866 532938 136102 533174
rect 136186 532938 136422 533174
rect 135866 497258 136102 497494
rect 136186 497258 136422 497494
rect 135866 496938 136102 497174
rect 136186 496938 136422 497174
rect 135866 461258 136102 461494
rect 136186 461258 136422 461494
rect 135866 460938 136102 461174
rect 136186 460938 136422 461174
rect 135866 425258 136102 425494
rect 136186 425258 136422 425494
rect 135866 424938 136102 425174
rect 136186 424938 136422 425174
rect 135866 389258 136102 389494
rect 136186 389258 136422 389494
rect 135866 388938 136102 389174
rect 136186 388938 136422 389174
rect 135866 353258 136102 353494
rect 136186 353258 136422 353494
rect 135866 352938 136102 353174
rect 136186 352938 136422 353174
rect 135866 317258 136102 317494
rect 136186 317258 136422 317494
rect 135866 316938 136102 317174
rect 136186 316938 136422 317174
rect 135866 281258 136102 281494
rect 136186 281258 136422 281494
rect 135866 280938 136102 281174
rect 136186 280938 136422 281174
rect 135866 245258 136102 245494
rect 136186 245258 136422 245494
rect 135866 244938 136102 245174
rect 136186 244938 136422 245174
rect 135866 209258 136102 209494
rect 136186 209258 136422 209494
rect 135866 208938 136102 209174
rect 136186 208938 136422 209174
rect 135866 173258 136102 173494
rect 136186 173258 136422 173494
rect 135866 172938 136102 173174
rect 136186 172938 136422 173174
rect 135866 137258 136102 137494
rect 136186 137258 136422 137494
rect 135866 136938 136102 137174
rect 136186 136938 136422 137174
rect 135866 101258 136102 101494
rect 136186 101258 136422 101494
rect 135866 100938 136102 101174
rect 136186 100938 136422 101174
rect 135866 65258 136102 65494
rect 136186 65258 136422 65494
rect 135866 64938 136102 65174
rect 136186 64938 136422 65174
rect 135866 29258 136102 29494
rect 136186 29258 136422 29494
rect 135866 28938 136102 29174
rect 136186 28938 136422 29174
rect 135866 -7302 136102 -7066
rect 136186 -7302 136422 -7066
rect 135866 -7622 136102 -7386
rect 136186 -7622 136422 -7386
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 705562 149782 705798
rect 149866 705562 150102 705798
rect 149546 705242 149782 705478
rect 149866 705242 150102 705478
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -1542 149782 -1306
rect 149866 -1542 150102 -1306
rect 149546 -1862 149782 -1626
rect 149866 -1862 150102 -1626
rect 153266 706522 153502 706758
rect 153586 706522 153822 706758
rect 153266 706202 153502 706438
rect 153586 706202 153822 706438
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -2502 153502 -2266
rect 153586 -2502 153822 -2266
rect 153266 -2822 153502 -2586
rect 153586 -2822 153822 -2586
rect 156986 707482 157222 707718
rect 157306 707482 157542 707718
rect 156986 707162 157222 707398
rect 157306 707162 157542 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 156986 -3462 157222 -3226
rect 157306 -3462 157542 -3226
rect 156986 -3782 157222 -3546
rect 157306 -3782 157542 -3546
rect 160706 708442 160942 708678
rect 161026 708442 161262 708678
rect 160706 708122 160942 708358
rect 161026 708122 161262 708358
rect 160706 666098 160942 666334
rect 161026 666098 161262 666334
rect 160706 665778 160942 666014
rect 161026 665778 161262 666014
rect 160706 630098 160942 630334
rect 161026 630098 161262 630334
rect 160706 629778 160942 630014
rect 161026 629778 161262 630014
rect 160706 594098 160942 594334
rect 161026 594098 161262 594334
rect 160706 593778 160942 594014
rect 161026 593778 161262 594014
rect 160706 558098 160942 558334
rect 161026 558098 161262 558334
rect 160706 557778 160942 558014
rect 161026 557778 161262 558014
rect 160706 522098 160942 522334
rect 161026 522098 161262 522334
rect 160706 521778 160942 522014
rect 161026 521778 161262 522014
rect 160706 486098 160942 486334
rect 161026 486098 161262 486334
rect 160706 485778 160942 486014
rect 161026 485778 161262 486014
rect 160706 450098 160942 450334
rect 161026 450098 161262 450334
rect 160706 449778 160942 450014
rect 161026 449778 161262 450014
rect 160706 414098 160942 414334
rect 161026 414098 161262 414334
rect 160706 413778 160942 414014
rect 161026 413778 161262 414014
rect 160706 378098 160942 378334
rect 161026 378098 161262 378334
rect 160706 377778 160942 378014
rect 161026 377778 161262 378014
rect 160706 342098 160942 342334
rect 161026 342098 161262 342334
rect 160706 341778 160942 342014
rect 161026 341778 161262 342014
rect 160706 306098 160942 306334
rect 161026 306098 161262 306334
rect 160706 305778 160942 306014
rect 161026 305778 161262 306014
rect 160706 270098 160942 270334
rect 161026 270098 161262 270334
rect 160706 269778 160942 270014
rect 161026 269778 161262 270014
rect 160706 234098 160942 234334
rect 161026 234098 161262 234334
rect 160706 233778 160942 234014
rect 161026 233778 161262 234014
rect 160706 198098 160942 198334
rect 161026 198098 161262 198334
rect 160706 197778 160942 198014
rect 161026 197778 161262 198014
rect 160706 162098 160942 162334
rect 161026 162098 161262 162334
rect 160706 161778 160942 162014
rect 161026 161778 161262 162014
rect 160706 126098 160942 126334
rect 161026 126098 161262 126334
rect 160706 125778 160942 126014
rect 161026 125778 161262 126014
rect 160706 90098 160942 90334
rect 161026 90098 161262 90334
rect 160706 89778 160942 90014
rect 161026 89778 161262 90014
rect 160706 54098 160942 54334
rect 161026 54098 161262 54334
rect 160706 53778 160942 54014
rect 161026 53778 161262 54014
rect 160706 18098 160942 18334
rect 161026 18098 161262 18334
rect 160706 17778 160942 18014
rect 161026 17778 161262 18014
rect 160706 -4422 160942 -4186
rect 161026 -4422 161262 -4186
rect 160706 -4742 160942 -4506
rect 161026 -4742 161262 -4506
rect 164426 709402 164662 709638
rect 164746 709402 164982 709638
rect 164426 709082 164662 709318
rect 164746 709082 164982 709318
rect 164426 669818 164662 670054
rect 164746 669818 164982 670054
rect 164426 669498 164662 669734
rect 164746 669498 164982 669734
rect 164426 633818 164662 634054
rect 164746 633818 164982 634054
rect 164426 633498 164662 633734
rect 164746 633498 164982 633734
rect 164426 597818 164662 598054
rect 164746 597818 164982 598054
rect 164426 597498 164662 597734
rect 164746 597498 164982 597734
rect 164426 561818 164662 562054
rect 164746 561818 164982 562054
rect 164426 561498 164662 561734
rect 164746 561498 164982 561734
rect 164426 525818 164662 526054
rect 164746 525818 164982 526054
rect 164426 525498 164662 525734
rect 164746 525498 164982 525734
rect 164426 489818 164662 490054
rect 164746 489818 164982 490054
rect 164426 489498 164662 489734
rect 164746 489498 164982 489734
rect 164426 453818 164662 454054
rect 164746 453818 164982 454054
rect 164426 453498 164662 453734
rect 164746 453498 164982 453734
rect 164426 417818 164662 418054
rect 164746 417818 164982 418054
rect 164426 417498 164662 417734
rect 164746 417498 164982 417734
rect 164426 381818 164662 382054
rect 164746 381818 164982 382054
rect 164426 381498 164662 381734
rect 164746 381498 164982 381734
rect 164426 345818 164662 346054
rect 164746 345818 164982 346054
rect 164426 345498 164662 345734
rect 164746 345498 164982 345734
rect 164426 309818 164662 310054
rect 164746 309818 164982 310054
rect 164426 309498 164662 309734
rect 164746 309498 164982 309734
rect 164426 273818 164662 274054
rect 164746 273818 164982 274054
rect 164426 273498 164662 273734
rect 164746 273498 164982 273734
rect 164426 237818 164662 238054
rect 164746 237818 164982 238054
rect 164426 237498 164662 237734
rect 164746 237498 164982 237734
rect 168146 710362 168382 710598
rect 168466 710362 168702 710598
rect 168146 710042 168382 710278
rect 168466 710042 168702 710278
rect 168146 673538 168382 673774
rect 168466 673538 168702 673774
rect 168146 673218 168382 673454
rect 168466 673218 168702 673454
rect 168146 637538 168382 637774
rect 168466 637538 168702 637774
rect 168146 637218 168382 637454
rect 168466 637218 168702 637454
rect 168146 601538 168382 601774
rect 168466 601538 168702 601774
rect 168146 601218 168382 601454
rect 168466 601218 168702 601454
rect 168146 565538 168382 565774
rect 168466 565538 168702 565774
rect 168146 565218 168382 565454
rect 168466 565218 168702 565454
rect 168146 529538 168382 529774
rect 168466 529538 168702 529774
rect 168146 529218 168382 529454
rect 168466 529218 168702 529454
rect 168146 493538 168382 493774
rect 168466 493538 168702 493774
rect 168146 493218 168382 493454
rect 168466 493218 168702 493454
rect 168146 457538 168382 457774
rect 168466 457538 168702 457774
rect 168146 457218 168382 457454
rect 168466 457218 168702 457454
rect 168146 421538 168382 421774
rect 168466 421538 168702 421774
rect 168146 421218 168382 421454
rect 168466 421218 168702 421454
rect 168146 385538 168382 385774
rect 168466 385538 168702 385774
rect 168146 385218 168382 385454
rect 168466 385218 168702 385454
rect 168146 349538 168382 349774
rect 168466 349538 168702 349774
rect 168146 349218 168382 349454
rect 168466 349218 168702 349454
rect 168146 313538 168382 313774
rect 168466 313538 168702 313774
rect 168146 313218 168382 313454
rect 168466 313218 168702 313454
rect 168146 277538 168382 277774
rect 168466 277538 168702 277774
rect 168146 277218 168382 277454
rect 168466 277218 168702 277454
rect 168146 241538 168382 241774
rect 168466 241538 168702 241774
rect 168146 241218 168382 241454
rect 168466 241218 168702 241454
rect 164426 201818 164662 202054
rect 164746 201818 164982 202054
rect 164426 201498 164662 201734
rect 164746 201498 164982 201734
rect 164426 165818 164662 166054
rect 164746 165818 164982 166054
rect 164426 165498 164662 165734
rect 164746 165498 164982 165734
rect 164426 129818 164662 130054
rect 164746 129818 164982 130054
rect 164426 129498 164662 129734
rect 164746 129498 164982 129734
rect 171866 711322 172102 711558
rect 172186 711322 172422 711558
rect 171866 711002 172102 711238
rect 172186 711002 172422 711238
rect 171866 677258 172102 677494
rect 172186 677258 172422 677494
rect 171866 676938 172102 677174
rect 172186 676938 172422 677174
rect 171866 641258 172102 641494
rect 172186 641258 172422 641494
rect 171866 640938 172102 641174
rect 172186 640938 172422 641174
rect 171866 605258 172102 605494
rect 172186 605258 172422 605494
rect 171866 604938 172102 605174
rect 172186 604938 172422 605174
rect 171866 569258 172102 569494
rect 172186 569258 172422 569494
rect 171866 568938 172102 569174
rect 172186 568938 172422 569174
rect 171866 533258 172102 533494
rect 172186 533258 172422 533494
rect 171866 532938 172102 533174
rect 172186 532938 172422 533174
rect 171866 497258 172102 497494
rect 172186 497258 172422 497494
rect 171866 496938 172102 497174
rect 172186 496938 172422 497174
rect 171866 461258 172102 461494
rect 172186 461258 172422 461494
rect 171866 460938 172102 461174
rect 172186 460938 172422 461174
rect 171866 425258 172102 425494
rect 172186 425258 172422 425494
rect 171866 424938 172102 425174
rect 172186 424938 172422 425174
rect 171866 389258 172102 389494
rect 172186 389258 172422 389494
rect 171866 388938 172102 389174
rect 172186 388938 172422 389174
rect 171866 353258 172102 353494
rect 172186 353258 172422 353494
rect 171866 352938 172102 353174
rect 172186 352938 172422 353174
rect 171866 317258 172102 317494
rect 172186 317258 172422 317494
rect 171866 316938 172102 317174
rect 172186 316938 172422 317174
rect 171866 281258 172102 281494
rect 172186 281258 172422 281494
rect 171866 280938 172102 281174
rect 172186 280938 172422 281174
rect 171866 245258 172102 245494
rect 172186 245258 172422 245494
rect 171866 244938 172102 245174
rect 172186 244938 172422 245174
rect 168146 205538 168382 205774
rect 168466 205538 168702 205774
rect 168146 205218 168382 205454
rect 168466 205218 168702 205454
rect 164426 93818 164662 94054
rect 164746 93818 164982 94054
rect 164426 93498 164662 93734
rect 164746 93498 164982 93734
rect 164426 57818 164662 58054
rect 164746 57818 164982 58054
rect 164426 57498 164662 57734
rect 164746 57498 164982 57734
rect 168146 169538 168382 169774
rect 168466 169538 168702 169774
rect 168146 169218 168382 169454
rect 168466 169218 168702 169454
rect 168146 133538 168382 133774
rect 168466 133538 168702 133774
rect 168146 133218 168382 133454
rect 168466 133218 168702 133454
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 174250 219218 174486 219454
rect 174250 218898 174486 219134
rect 185546 705562 185782 705798
rect 185866 705562 186102 705798
rect 185546 705242 185782 705478
rect 185866 705242 186102 705478
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 189266 706522 189502 706758
rect 189586 706522 189822 706758
rect 189266 706202 189502 706438
rect 189586 706202 189822 706438
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 192986 707482 193222 707718
rect 193306 707482 193542 707718
rect 192986 707162 193222 707398
rect 193306 707162 193542 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 196706 708442 196942 708678
rect 197026 708442 197262 708678
rect 196706 708122 196942 708358
rect 197026 708122 197262 708358
rect 196706 666098 196942 666334
rect 197026 666098 197262 666334
rect 196706 665778 196942 666014
rect 197026 665778 197262 666014
rect 196706 630098 196942 630334
rect 197026 630098 197262 630334
rect 196706 629778 196942 630014
rect 197026 629778 197262 630014
rect 196706 594098 196942 594334
rect 197026 594098 197262 594334
rect 196706 593778 196942 594014
rect 197026 593778 197262 594014
rect 196706 558098 196942 558334
rect 197026 558098 197262 558334
rect 196706 557778 196942 558014
rect 197026 557778 197262 558014
rect 196706 522098 196942 522334
rect 197026 522098 197262 522334
rect 196706 521778 196942 522014
rect 197026 521778 197262 522014
rect 196706 486098 196942 486334
rect 197026 486098 197262 486334
rect 196706 485778 196942 486014
rect 197026 485778 197262 486014
rect 196706 450098 196942 450334
rect 197026 450098 197262 450334
rect 196706 449778 196942 450014
rect 197026 449778 197262 450014
rect 196706 414098 196942 414334
rect 197026 414098 197262 414334
rect 196706 413778 196942 414014
rect 197026 413778 197262 414014
rect 196706 378098 196942 378334
rect 197026 378098 197262 378334
rect 196706 377778 196942 378014
rect 197026 377778 197262 378014
rect 196706 342098 196942 342334
rect 197026 342098 197262 342334
rect 196706 341778 196942 342014
rect 197026 341778 197262 342014
rect 196706 306098 196942 306334
rect 197026 306098 197262 306334
rect 196706 305778 196942 306014
rect 197026 305778 197262 306014
rect 196706 270098 196942 270334
rect 197026 270098 197262 270334
rect 196706 269778 196942 270014
rect 197026 269778 197262 270014
rect 196706 234098 196942 234334
rect 197026 234098 197262 234334
rect 196706 233778 196942 234014
rect 197026 233778 197262 234014
rect 200426 709402 200662 709638
rect 200746 709402 200982 709638
rect 200426 709082 200662 709318
rect 200746 709082 200982 709318
rect 200426 669818 200662 670054
rect 200746 669818 200982 670054
rect 200426 669498 200662 669734
rect 200746 669498 200982 669734
rect 200426 633818 200662 634054
rect 200746 633818 200982 634054
rect 200426 633498 200662 633734
rect 200746 633498 200982 633734
rect 200426 597818 200662 598054
rect 200746 597818 200982 598054
rect 200426 597498 200662 597734
rect 200746 597498 200982 597734
rect 200426 561818 200662 562054
rect 200746 561818 200982 562054
rect 200426 561498 200662 561734
rect 200746 561498 200982 561734
rect 200426 525818 200662 526054
rect 200746 525818 200982 526054
rect 200426 525498 200662 525734
rect 200746 525498 200982 525734
rect 200426 489818 200662 490054
rect 200746 489818 200982 490054
rect 200426 489498 200662 489734
rect 200746 489498 200982 489734
rect 200426 453818 200662 454054
rect 200746 453818 200982 454054
rect 200426 453498 200662 453734
rect 200746 453498 200982 453734
rect 200426 417818 200662 418054
rect 200746 417818 200982 418054
rect 200426 417498 200662 417734
rect 200746 417498 200982 417734
rect 200426 381818 200662 382054
rect 200746 381818 200982 382054
rect 200426 381498 200662 381734
rect 200746 381498 200982 381734
rect 200426 345818 200662 346054
rect 200746 345818 200982 346054
rect 200426 345498 200662 345734
rect 200746 345498 200982 345734
rect 200426 309818 200662 310054
rect 200746 309818 200982 310054
rect 200426 309498 200662 309734
rect 200746 309498 200982 309734
rect 200426 273818 200662 274054
rect 200746 273818 200982 274054
rect 200426 273498 200662 273734
rect 200746 273498 200982 273734
rect 200426 237818 200662 238054
rect 200746 237818 200982 238054
rect 200426 237498 200662 237734
rect 200746 237498 200982 237734
rect 204146 710362 204382 710598
rect 204466 710362 204702 710598
rect 204146 710042 204382 710278
rect 204466 710042 204702 710278
rect 204146 673538 204382 673774
rect 204466 673538 204702 673774
rect 204146 673218 204382 673454
rect 204466 673218 204702 673454
rect 204146 637538 204382 637774
rect 204466 637538 204702 637774
rect 204146 637218 204382 637454
rect 204466 637218 204702 637454
rect 204146 601538 204382 601774
rect 204466 601538 204702 601774
rect 204146 601218 204382 601454
rect 204466 601218 204702 601454
rect 204146 565538 204382 565774
rect 204466 565538 204702 565774
rect 204146 565218 204382 565454
rect 204466 565218 204702 565454
rect 204146 529538 204382 529774
rect 204466 529538 204702 529774
rect 204146 529218 204382 529454
rect 204466 529218 204702 529454
rect 204146 493538 204382 493774
rect 204466 493538 204702 493774
rect 204146 493218 204382 493454
rect 204466 493218 204702 493454
rect 204146 457538 204382 457774
rect 204466 457538 204702 457774
rect 204146 457218 204382 457454
rect 204466 457218 204702 457454
rect 204146 421538 204382 421774
rect 204466 421538 204702 421774
rect 204146 421218 204382 421454
rect 204466 421218 204702 421454
rect 204146 385538 204382 385774
rect 204466 385538 204702 385774
rect 204146 385218 204382 385454
rect 204466 385218 204702 385454
rect 204146 349538 204382 349774
rect 204466 349538 204702 349774
rect 204146 349218 204382 349454
rect 204466 349218 204702 349454
rect 204146 313538 204382 313774
rect 204466 313538 204702 313774
rect 204146 313218 204382 313454
rect 204466 313218 204702 313454
rect 204146 277538 204382 277774
rect 204466 277538 204702 277774
rect 204146 277218 204382 277454
rect 204466 277218 204702 277454
rect 204146 241538 204382 241774
rect 204466 241538 204702 241774
rect 204146 241218 204382 241454
rect 204466 241218 204702 241454
rect 207866 711322 208102 711558
rect 208186 711322 208422 711558
rect 207866 711002 208102 711238
rect 208186 711002 208422 711238
rect 207866 677258 208102 677494
rect 208186 677258 208422 677494
rect 207866 676938 208102 677174
rect 208186 676938 208422 677174
rect 207866 641258 208102 641494
rect 208186 641258 208422 641494
rect 207866 640938 208102 641174
rect 208186 640938 208422 641174
rect 207866 605258 208102 605494
rect 208186 605258 208422 605494
rect 207866 604938 208102 605174
rect 208186 604938 208422 605174
rect 207866 569258 208102 569494
rect 208186 569258 208422 569494
rect 207866 568938 208102 569174
rect 208186 568938 208422 569174
rect 207866 533258 208102 533494
rect 208186 533258 208422 533494
rect 207866 532938 208102 533174
rect 208186 532938 208422 533174
rect 207866 497258 208102 497494
rect 208186 497258 208422 497494
rect 207866 496938 208102 497174
rect 208186 496938 208422 497174
rect 207866 461258 208102 461494
rect 208186 461258 208422 461494
rect 207866 460938 208102 461174
rect 208186 460938 208422 461174
rect 207866 425258 208102 425494
rect 208186 425258 208422 425494
rect 207866 424938 208102 425174
rect 208186 424938 208422 425174
rect 207866 389258 208102 389494
rect 208186 389258 208422 389494
rect 207866 388938 208102 389174
rect 208186 388938 208422 389174
rect 207866 353258 208102 353494
rect 208186 353258 208422 353494
rect 207866 352938 208102 353174
rect 208186 352938 208422 353174
rect 207866 317258 208102 317494
rect 208186 317258 208422 317494
rect 207866 316938 208102 317174
rect 208186 316938 208422 317174
rect 207866 281258 208102 281494
rect 208186 281258 208422 281494
rect 207866 280938 208102 281174
rect 208186 280938 208422 281174
rect 207866 245258 208102 245494
rect 208186 245258 208422 245494
rect 207866 244938 208102 245174
rect 208186 244938 208422 245174
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 221546 705562 221782 705798
rect 221866 705562 222102 705798
rect 221546 705242 221782 705478
rect 221866 705242 222102 705478
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 189610 222938 189846 223174
rect 189610 222618 189846 222854
rect 220330 222938 220566 223174
rect 220330 222618 220566 222854
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 171866 209258 172102 209494
rect 172186 209258 172422 209494
rect 171866 208938 172102 209174
rect 172186 208938 172422 209174
rect 174250 183218 174486 183454
rect 174250 182898 174486 183134
rect 204970 219218 205206 219454
rect 204970 218898 205206 219134
rect 189610 186938 189846 187174
rect 189610 186618 189846 186854
rect 220330 186938 220566 187174
rect 220330 186618 220566 186854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 171866 173258 172102 173494
rect 172186 173258 172422 173494
rect 171866 172938 172102 173174
rect 172186 172938 172422 173174
rect 171866 137258 172102 137494
rect 172186 137258 172422 137494
rect 171866 136938 172102 137174
rect 172186 136938 172422 137174
rect 168146 97538 168382 97774
rect 168466 97538 168702 97774
rect 168146 97218 168382 97454
rect 168466 97218 168702 97454
rect 168146 61538 168382 61774
rect 168466 61538 168702 61774
rect 168146 61218 168382 61454
rect 168466 61218 168702 61454
rect 164426 21818 164662 22054
rect 164746 21818 164982 22054
rect 164426 21498 164662 21734
rect 164746 21498 164982 21734
rect 164426 -5382 164662 -5146
rect 164746 -5382 164982 -5146
rect 164426 -5702 164662 -5466
rect 164746 -5702 164982 -5466
rect 168146 25538 168382 25774
rect 168466 25538 168702 25774
rect 168146 25218 168382 25454
rect 168466 25218 168702 25454
rect 204970 183218 205206 183454
rect 204970 182898 205206 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 177932 114938 178168 115174
rect 177932 114618 178168 114854
rect 174459 111218 174695 111454
rect 174459 110898 174695 111134
rect 181405 111218 181641 111454
rect 181405 110898 181641 111134
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 184878 114938 185114 115174
rect 184878 114618 185114 114854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 171866 101258 172102 101494
rect 172186 101258 172422 101494
rect 171866 100938 172102 101174
rect 172186 100938 172422 101174
rect 177932 78938 178168 79174
rect 177932 78618 178168 78854
rect 174459 75218 174695 75454
rect 174459 74898 174695 75134
rect 181405 75218 181641 75454
rect 181405 74898 181641 75134
rect 184878 78938 185114 79174
rect 184878 78618 185114 78854
rect 191824 114938 192060 115174
rect 191824 114618 192060 114854
rect 188351 111218 188587 111454
rect 188351 110898 188587 111134
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 171866 65258 172102 65494
rect 172186 65258 172422 65494
rect 171866 64938 172102 65174
rect 172186 64938 172422 65174
rect 171866 29258 172102 29494
rect 172186 29258 172422 29494
rect 171866 28938 172102 29174
rect 172186 28938 172422 29174
rect 168146 -6342 168382 -6106
rect 168466 -6342 168702 -6106
rect 168146 -6662 168382 -6426
rect 168466 -6662 168702 -6426
rect 171866 -7302 172102 -7066
rect 172186 -7302 172422 -7066
rect 171866 -7622 172102 -7386
rect 172186 -7622 172422 -7386
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 188351 75218 188587 75454
rect 188351 74898 188587 75134
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -1542 185782 -1306
rect 185866 -1542 186102 -1306
rect 185546 -1862 185782 -1626
rect 185866 -1862 186102 -1626
rect 196706 162098 196942 162334
rect 197026 162098 197262 162334
rect 196706 161778 196942 162014
rect 197026 161778 197262 162014
rect 196706 126098 196942 126334
rect 197026 126098 197262 126334
rect 196706 125778 196942 126014
rect 197026 125778 197262 126014
rect 195297 111218 195533 111454
rect 195297 110898 195533 111134
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 191824 78938 192060 79174
rect 191824 78618 192060 78854
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -2502 189502 -2266
rect 189586 -2502 189822 -2266
rect 189266 -2822 189502 -2586
rect 189586 -2822 189822 -2586
rect 198770 114938 199006 115174
rect 198770 114618 199006 114854
rect 200426 165818 200662 166054
rect 200746 165818 200982 166054
rect 200426 165498 200662 165734
rect 200746 165498 200982 165734
rect 200426 129818 200662 130054
rect 200746 129818 200982 130054
rect 200426 129498 200662 129734
rect 200746 129498 200982 129734
rect 204146 169538 204382 169774
rect 204466 169538 204702 169774
rect 204146 169218 204382 169454
rect 204466 169218 204702 169454
rect 204146 133538 204382 133774
rect 204466 133538 204702 133774
rect 204146 133218 204382 133454
rect 204466 133218 204702 133454
rect 200426 93818 200662 94054
rect 200746 93818 200982 94054
rect 200426 93498 200662 93734
rect 200746 93498 200982 93734
rect 196706 90098 196942 90334
rect 197026 90098 197262 90334
rect 196706 89778 196942 90014
rect 197026 89778 197262 90014
rect 195297 75218 195533 75454
rect 195297 74898 195533 75134
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 192986 -3462 193222 -3226
rect 193306 -3462 193542 -3226
rect 192986 -3782 193222 -3546
rect 193306 -3782 193542 -3546
rect 198770 78938 199006 79174
rect 198770 78618 199006 78854
rect 196706 54098 196942 54334
rect 197026 54098 197262 54334
rect 196706 53778 196942 54014
rect 197026 53778 197262 54014
rect 196706 18098 196942 18334
rect 197026 18098 197262 18334
rect 196706 17778 196942 18014
rect 197026 17778 197262 18014
rect 196706 -4422 196942 -4186
rect 197026 -4422 197262 -4186
rect 196706 -4742 196942 -4506
rect 197026 -4742 197262 -4506
rect 204146 97538 204382 97774
rect 204466 97538 204702 97774
rect 204146 97218 204382 97454
rect 204466 97218 204702 97454
rect 200426 57818 200662 58054
rect 200746 57818 200982 58054
rect 200426 57498 200662 57734
rect 200746 57498 200982 57734
rect 200426 21818 200662 22054
rect 200746 21818 200982 22054
rect 200426 21498 200662 21734
rect 200746 21498 200982 21734
rect 200426 -5382 200662 -5146
rect 200746 -5382 200982 -5146
rect 200426 -5702 200662 -5466
rect 200746 -5702 200982 -5466
rect 204146 61538 204382 61774
rect 204466 61538 204702 61774
rect 204146 61218 204382 61454
rect 204466 61218 204702 61454
rect 204146 25538 204382 25774
rect 204466 25538 204702 25774
rect 204146 25218 204382 25454
rect 204466 25218 204702 25454
rect 204146 -6342 204382 -6106
rect 204466 -6342 204702 -6106
rect 204146 -6662 204382 -6426
rect 204466 -6662 204702 -6426
rect 207866 173258 208102 173494
rect 208186 173258 208422 173494
rect 207866 172938 208102 173174
rect 208186 172938 208422 173174
rect 207866 137258 208102 137494
rect 208186 137258 208422 137494
rect 207866 136938 208102 137174
rect 208186 136938 208422 137174
rect 207866 101258 208102 101494
rect 208186 101258 208422 101494
rect 207866 100938 208102 101174
rect 208186 100938 208422 101174
rect 207866 65258 208102 65494
rect 208186 65258 208422 65494
rect 207866 64938 208102 65174
rect 208186 64938 208422 65174
rect 207866 29258 208102 29494
rect 208186 29258 208422 29494
rect 207866 28938 208102 29174
rect 208186 28938 208422 29174
rect 207866 -7302 208102 -7066
rect 208186 -7302 208422 -7066
rect 207866 -7622 208102 -7386
rect 208186 -7622 208422 -7386
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -1542 221782 -1306
rect 221866 -1542 222102 -1306
rect 221546 -1862 221782 -1626
rect 221866 -1862 222102 -1626
rect 225266 706522 225502 706758
rect 225586 706522 225822 706758
rect 225266 706202 225502 706438
rect 225586 706202 225822 706438
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 225266 118658 225502 118894
rect 225586 118658 225822 118894
rect 225266 118338 225502 118574
rect 225586 118338 225822 118574
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -2502 225502 -2266
rect 225586 -2502 225822 -2266
rect 225266 -2822 225502 -2586
rect 225586 -2822 225822 -2586
rect 228986 707482 229222 707718
rect 229306 707482 229542 707718
rect 228986 707162 229222 707398
rect 229306 707162 229542 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 232706 708442 232942 708678
rect 233026 708442 233262 708678
rect 232706 708122 232942 708358
rect 233026 708122 233262 708358
rect 232706 666098 232942 666334
rect 233026 666098 233262 666334
rect 232706 665778 232942 666014
rect 233026 665778 233262 666014
rect 232706 630098 232942 630334
rect 233026 630098 233262 630334
rect 232706 629778 232942 630014
rect 233026 629778 233262 630014
rect 232706 594098 232942 594334
rect 233026 594098 233262 594334
rect 232706 593778 232942 594014
rect 233026 593778 233262 594014
rect 232706 558098 232942 558334
rect 233026 558098 233262 558334
rect 232706 557778 232942 558014
rect 233026 557778 233262 558014
rect 232706 522098 232942 522334
rect 233026 522098 233262 522334
rect 232706 521778 232942 522014
rect 233026 521778 233262 522014
rect 232706 486098 232942 486334
rect 233026 486098 233262 486334
rect 232706 485778 232942 486014
rect 233026 485778 233262 486014
rect 232706 450098 232942 450334
rect 233026 450098 233262 450334
rect 232706 449778 232942 450014
rect 233026 449778 233262 450014
rect 232706 414098 232942 414334
rect 233026 414098 233262 414334
rect 232706 413778 232942 414014
rect 233026 413778 233262 414014
rect 232706 378098 232942 378334
rect 233026 378098 233262 378334
rect 232706 377778 232942 378014
rect 233026 377778 233262 378014
rect 232706 342098 232942 342334
rect 233026 342098 233262 342334
rect 232706 341778 232942 342014
rect 233026 341778 233262 342014
rect 232706 306098 232942 306334
rect 233026 306098 233262 306334
rect 232706 305778 232942 306014
rect 233026 305778 233262 306014
rect 232706 270098 232942 270334
rect 233026 270098 233262 270334
rect 232706 269778 232942 270014
rect 233026 269778 233262 270014
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 232706 234098 232942 234334
rect 233026 234098 233262 234334
rect 232706 233778 232942 234014
rect 233026 233778 233262 234014
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 228986 -3462 229222 -3226
rect 229306 -3462 229542 -3226
rect 228986 -3782 229222 -3546
rect 229306 -3782 229542 -3546
rect 232706 198098 232942 198334
rect 233026 198098 233262 198334
rect 232706 197778 232942 198014
rect 233026 197778 233262 198014
rect 232706 162098 232942 162334
rect 233026 162098 233262 162334
rect 232706 161778 232942 162014
rect 233026 161778 233262 162014
rect 232706 126098 232942 126334
rect 233026 126098 233262 126334
rect 232706 125778 232942 126014
rect 233026 125778 233262 126014
rect 232706 90098 232942 90334
rect 233026 90098 233262 90334
rect 232706 89778 232942 90014
rect 233026 89778 233262 90014
rect 232706 54098 232942 54334
rect 233026 54098 233262 54334
rect 232706 53778 232942 54014
rect 233026 53778 233262 54014
rect 232706 18098 232942 18334
rect 233026 18098 233262 18334
rect 232706 17778 232942 18014
rect 233026 17778 233262 18014
rect 232706 -4422 232942 -4186
rect 233026 -4422 233262 -4186
rect 232706 -4742 232942 -4506
rect 233026 -4742 233262 -4506
rect 236426 709402 236662 709638
rect 236746 709402 236982 709638
rect 236426 709082 236662 709318
rect 236746 709082 236982 709318
rect 236426 669818 236662 670054
rect 236746 669818 236982 670054
rect 236426 669498 236662 669734
rect 236746 669498 236982 669734
rect 236426 633818 236662 634054
rect 236746 633818 236982 634054
rect 236426 633498 236662 633734
rect 236746 633498 236982 633734
rect 236426 597818 236662 598054
rect 236746 597818 236982 598054
rect 236426 597498 236662 597734
rect 236746 597498 236982 597734
rect 236426 561818 236662 562054
rect 236746 561818 236982 562054
rect 236426 561498 236662 561734
rect 236746 561498 236982 561734
rect 236426 525818 236662 526054
rect 236746 525818 236982 526054
rect 236426 525498 236662 525734
rect 236746 525498 236982 525734
rect 236426 489818 236662 490054
rect 236746 489818 236982 490054
rect 236426 489498 236662 489734
rect 236746 489498 236982 489734
rect 236426 453818 236662 454054
rect 236746 453818 236982 454054
rect 236426 453498 236662 453734
rect 236746 453498 236982 453734
rect 236426 417818 236662 418054
rect 236746 417818 236982 418054
rect 236426 417498 236662 417734
rect 236746 417498 236982 417734
rect 236426 381818 236662 382054
rect 236746 381818 236982 382054
rect 236426 381498 236662 381734
rect 236746 381498 236982 381734
rect 236426 345818 236662 346054
rect 236746 345818 236982 346054
rect 236426 345498 236662 345734
rect 236746 345498 236982 345734
rect 236426 309818 236662 310054
rect 236746 309818 236982 310054
rect 236426 309498 236662 309734
rect 236746 309498 236982 309734
rect 236426 273818 236662 274054
rect 236746 273818 236982 274054
rect 236426 273498 236662 273734
rect 236746 273498 236982 273734
rect 236426 237818 236662 238054
rect 236746 237818 236982 238054
rect 236426 237498 236662 237734
rect 236746 237498 236982 237734
rect 236426 201818 236662 202054
rect 236746 201818 236982 202054
rect 236426 201498 236662 201734
rect 236746 201498 236982 201734
rect 236426 165818 236662 166054
rect 236746 165818 236982 166054
rect 236426 165498 236662 165734
rect 236746 165498 236982 165734
rect 236426 129818 236662 130054
rect 236746 129818 236982 130054
rect 236426 129498 236662 129734
rect 236746 129498 236982 129734
rect 236426 93818 236662 94054
rect 236746 93818 236982 94054
rect 236426 93498 236662 93734
rect 236746 93498 236982 93734
rect 236426 57818 236662 58054
rect 236746 57818 236982 58054
rect 236426 57498 236662 57734
rect 236746 57498 236982 57734
rect 236426 21818 236662 22054
rect 236746 21818 236982 22054
rect 236426 21498 236662 21734
rect 236746 21498 236982 21734
rect 236426 -5382 236662 -5146
rect 236746 -5382 236982 -5146
rect 236426 -5702 236662 -5466
rect 236746 -5702 236982 -5466
rect 240146 710362 240382 710598
rect 240466 710362 240702 710598
rect 240146 710042 240382 710278
rect 240466 710042 240702 710278
rect 240146 673538 240382 673774
rect 240466 673538 240702 673774
rect 240146 673218 240382 673454
rect 240466 673218 240702 673454
rect 240146 637538 240382 637774
rect 240466 637538 240702 637774
rect 240146 637218 240382 637454
rect 240466 637218 240702 637454
rect 240146 601538 240382 601774
rect 240466 601538 240702 601774
rect 240146 601218 240382 601454
rect 240466 601218 240702 601454
rect 240146 565538 240382 565774
rect 240466 565538 240702 565774
rect 240146 565218 240382 565454
rect 240466 565218 240702 565454
rect 240146 529538 240382 529774
rect 240466 529538 240702 529774
rect 240146 529218 240382 529454
rect 240466 529218 240702 529454
rect 240146 493538 240382 493774
rect 240466 493538 240702 493774
rect 240146 493218 240382 493454
rect 240466 493218 240702 493454
rect 240146 457538 240382 457774
rect 240466 457538 240702 457774
rect 240146 457218 240382 457454
rect 240466 457218 240702 457454
rect 240146 421538 240382 421774
rect 240466 421538 240702 421774
rect 240146 421218 240382 421454
rect 240466 421218 240702 421454
rect 240146 385538 240382 385774
rect 240466 385538 240702 385774
rect 240146 385218 240382 385454
rect 240466 385218 240702 385454
rect 240146 349538 240382 349774
rect 240466 349538 240702 349774
rect 240146 349218 240382 349454
rect 240466 349218 240702 349454
rect 240146 313538 240382 313774
rect 240466 313538 240702 313774
rect 240146 313218 240382 313454
rect 240466 313218 240702 313454
rect 240146 277538 240382 277774
rect 240466 277538 240702 277774
rect 240146 277218 240382 277454
rect 240466 277218 240702 277454
rect 240146 241538 240382 241774
rect 240466 241538 240702 241774
rect 240146 241218 240382 241454
rect 240466 241218 240702 241454
rect 240146 205538 240382 205774
rect 240466 205538 240702 205774
rect 240146 205218 240382 205454
rect 240466 205218 240702 205454
rect 240146 169538 240382 169774
rect 240466 169538 240702 169774
rect 240146 169218 240382 169454
rect 240466 169218 240702 169454
rect 240146 133538 240382 133774
rect 240466 133538 240702 133774
rect 240146 133218 240382 133454
rect 240466 133218 240702 133454
rect 240146 97538 240382 97774
rect 240466 97538 240702 97774
rect 240146 97218 240382 97454
rect 240466 97218 240702 97454
rect 240146 61538 240382 61774
rect 240466 61538 240702 61774
rect 240146 61218 240382 61454
rect 240466 61218 240702 61454
rect 240146 25538 240382 25774
rect 240466 25538 240702 25774
rect 240146 25218 240382 25454
rect 240466 25218 240702 25454
rect 240146 -6342 240382 -6106
rect 240466 -6342 240702 -6106
rect 240146 -6662 240382 -6426
rect 240466 -6662 240702 -6426
rect 243866 711322 244102 711558
rect 244186 711322 244422 711558
rect 243866 711002 244102 711238
rect 244186 711002 244422 711238
rect 243866 677258 244102 677494
rect 244186 677258 244422 677494
rect 243866 676938 244102 677174
rect 244186 676938 244422 677174
rect 243866 641258 244102 641494
rect 244186 641258 244422 641494
rect 243866 640938 244102 641174
rect 244186 640938 244422 641174
rect 243866 605258 244102 605494
rect 244186 605258 244422 605494
rect 243866 604938 244102 605174
rect 244186 604938 244422 605174
rect 243866 569258 244102 569494
rect 244186 569258 244422 569494
rect 243866 568938 244102 569174
rect 244186 568938 244422 569174
rect 243866 533258 244102 533494
rect 244186 533258 244422 533494
rect 243866 532938 244102 533174
rect 244186 532938 244422 533174
rect 243866 497258 244102 497494
rect 244186 497258 244422 497494
rect 243866 496938 244102 497174
rect 244186 496938 244422 497174
rect 243866 461258 244102 461494
rect 244186 461258 244422 461494
rect 243866 460938 244102 461174
rect 244186 460938 244422 461174
rect 243866 425258 244102 425494
rect 244186 425258 244422 425494
rect 243866 424938 244102 425174
rect 244186 424938 244422 425174
rect 243866 389258 244102 389494
rect 244186 389258 244422 389494
rect 243866 388938 244102 389174
rect 244186 388938 244422 389174
rect 243866 353258 244102 353494
rect 244186 353258 244422 353494
rect 243866 352938 244102 353174
rect 244186 352938 244422 353174
rect 243866 317258 244102 317494
rect 244186 317258 244422 317494
rect 243866 316938 244102 317174
rect 244186 316938 244422 317174
rect 243866 281258 244102 281494
rect 244186 281258 244422 281494
rect 243866 280938 244102 281174
rect 244186 280938 244422 281174
rect 243866 245258 244102 245494
rect 244186 245258 244422 245494
rect 243866 244938 244102 245174
rect 244186 244938 244422 245174
rect 243866 209258 244102 209494
rect 244186 209258 244422 209494
rect 243866 208938 244102 209174
rect 244186 208938 244422 209174
rect 243866 173258 244102 173494
rect 244186 173258 244422 173494
rect 243866 172938 244102 173174
rect 244186 172938 244422 173174
rect 243866 137258 244102 137494
rect 244186 137258 244422 137494
rect 243866 136938 244102 137174
rect 244186 136938 244422 137174
rect 243866 101258 244102 101494
rect 244186 101258 244422 101494
rect 243866 100938 244102 101174
rect 244186 100938 244422 101174
rect 243866 65258 244102 65494
rect 244186 65258 244422 65494
rect 243866 64938 244102 65174
rect 244186 64938 244422 65174
rect 243866 29258 244102 29494
rect 244186 29258 244422 29494
rect 243866 28938 244102 29174
rect 244186 28938 244422 29174
rect 243866 -7302 244102 -7066
rect 244186 -7302 244422 -7066
rect 243866 -7622 244102 -7386
rect 244186 -7622 244422 -7386
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 705562 257782 705798
rect 257866 705562 258102 705798
rect 257546 705242 257782 705478
rect 257866 705242 258102 705478
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -1542 257782 -1306
rect 257866 -1542 258102 -1306
rect 257546 -1862 257782 -1626
rect 257866 -1862 258102 -1626
rect 261266 706522 261502 706758
rect 261586 706522 261822 706758
rect 261266 706202 261502 706438
rect 261586 706202 261822 706438
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -2502 261502 -2266
rect 261586 -2502 261822 -2266
rect 261266 -2822 261502 -2586
rect 261586 -2822 261822 -2586
rect 264986 707482 265222 707718
rect 265306 707482 265542 707718
rect 264986 707162 265222 707398
rect 265306 707162 265542 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 264986 -3462 265222 -3226
rect 265306 -3462 265542 -3226
rect 264986 -3782 265222 -3546
rect 265306 -3782 265542 -3546
rect 268706 708442 268942 708678
rect 269026 708442 269262 708678
rect 268706 708122 268942 708358
rect 269026 708122 269262 708358
rect 268706 666098 268942 666334
rect 269026 666098 269262 666334
rect 268706 665778 268942 666014
rect 269026 665778 269262 666014
rect 268706 630098 268942 630334
rect 269026 630098 269262 630334
rect 268706 629778 268942 630014
rect 269026 629778 269262 630014
rect 268706 594098 268942 594334
rect 269026 594098 269262 594334
rect 268706 593778 268942 594014
rect 269026 593778 269262 594014
rect 268706 558098 268942 558334
rect 269026 558098 269262 558334
rect 268706 557778 268942 558014
rect 269026 557778 269262 558014
rect 268706 522098 268942 522334
rect 269026 522098 269262 522334
rect 268706 521778 268942 522014
rect 269026 521778 269262 522014
rect 268706 486098 268942 486334
rect 269026 486098 269262 486334
rect 268706 485778 268942 486014
rect 269026 485778 269262 486014
rect 268706 450098 268942 450334
rect 269026 450098 269262 450334
rect 268706 449778 268942 450014
rect 269026 449778 269262 450014
rect 268706 414098 268942 414334
rect 269026 414098 269262 414334
rect 268706 413778 268942 414014
rect 269026 413778 269262 414014
rect 268706 378098 268942 378334
rect 269026 378098 269262 378334
rect 268706 377778 268942 378014
rect 269026 377778 269262 378014
rect 268706 342098 268942 342334
rect 269026 342098 269262 342334
rect 268706 341778 268942 342014
rect 269026 341778 269262 342014
rect 268706 306098 268942 306334
rect 269026 306098 269262 306334
rect 268706 305778 268942 306014
rect 269026 305778 269262 306014
rect 268706 270098 268942 270334
rect 269026 270098 269262 270334
rect 268706 269778 268942 270014
rect 269026 269778 269262 270014
rect 268706 234098 268942 234334
rect 269026 234098 269262 234334
rect 268706 233778 268942 234014
rect 269026 233778 269262 234014
rect 268706 198098 268942 198334
rect 269026 198098 269262 198334
rect 268706 197778 268942 198014
rect 269026 197778 269262 198014
rect 268706 162098 268942 162334
rect 269026 162098 269262 162334
rect 268706 161778 268942 162014
rect 269026 161778 269262 162014
rect 268706 126098 268942 126334
rect 269026 126098 269262 126334
rect 268706 125778 268942 126014
rect 269026 125778 269262 126014
rect 268706 90098 268942 90334
rect 269026 90098 269262 90334
rect 268706 89778 268942 90014
rect 269026 89778 269262 90014
rect 268706 54098 268942 54334
rect 269026 54098 269262 54334
rect 268706 53778 268942 54014
rect 269026 53778 269262 54014
rect 268706 18098 268942 18334
rect 269026 18098 269262 18334
rect 268706 17778 268942 18014
rect 269026 17778 269262 18014
rect 268706 -4422 268942 -4186
rect 269026 -4422 269262 -4186
rect 268706 -4742 268942 -4506
rect 269026 -4742 269262 -4506
rect 272426 709402 272662 709638
rect 272746 709402 272982 709638
rect 272426 709082 272662 709318
rect 272746 709082 272982 709318
rect 272426 669818 272662 670054
rect 272746 669818 272982 670054
rect 272426 669498 272662 669734
rect 272746 669498 272982 669734
rect 272426 633818 272662 634054
rect 272746 633818 272982 634054
rect 272426 633498 272662 633734
rect 272746 633498 272982 633734
rect 272426 597818 272662 598054
rect 272746 597818 272982 598054
rect 272426 597498 272662 597734
rect 272746 597498 272982 597734
rect 272426 561818 272662 562054
rect 272746 561818 272982 562054
rect 272426 561498 272662 561734
rect 272746 561498 272982 561734
rect 272426 525818 272662 526054
rect 272746 525818 272982 526054
rect 272426 525498 272662 525734
rect 272746 525498 272982 525734
rect 272426 489818 272662 490054
rect 272746 489818 272982 490054
rect 272426 489498 272662 489734
rect 272746 489498 272982 489734
rect 272426 453818 272662 454054
rect 272746 453818 272982 454054
rect 272426 453498 272662 453734
rect 272746 453498 272982 453734
rect 272426 417818 272662 418054
rect 272746 417818 272982 418054
rect 272426 417498 272662 417734
rect 272746 417498 272982 417734
rect 272426 381818 272662 382054
rect 272746 381818 272982 382054
rect 272426 381498 272662 381734
rect 272746 381498 272982 381734
rect 272426 345818 272662 346054
rect 272746 345818 272982 346054
rect 272426 345498 272662 345734
rect 272746 345498 272982 345734
rect 272426 309818 272662 310054
rect 272746 309818 272982 310054
rect 272426 309498 272662 309734
rect 272746 309498 272982 309734
rect 272426 273818 272662 274054
rect 272746 273818 272982 274054
rect 272426 273498 272662 273734
rect 272746 273498 272982 273734
rect 272426 237818 272662 238054
rect 272746 237818 272982 238054
rect 272426 237498 272662 237734
rect 272746 237498 272982 237734
rect 272426 201818 272662 202054
rect 272746 201818 272982 202054
rect 272426 201498 272662 201734
rect 272746 201498 272982 201734
rect 272426 165818 272662 166054
rect 272746 165818 272982 166054
rect 272426 165498 272662 165734
rect 272746 165498 272982 165734
rect 272426 129818 272662 130054
rect 272746 129818 272982 130054
rect 272426 129498 272662 129734
rect 272746 129498 272982 129734
rect 272426 93818 272662 94054
rect 272746 93818 272982 94054
rect 272426 93498 272662 93734
rect 272746 93498 272982 93734
rect 272426 57818 272662 58054
rect 272746 57818 272982 58054
rect 272426 57498 272662 57734
rect 272746 57498 272982 57734
rect 272426 21818 272662 22054
rect 272746 21818 272982 22054
rect 272426 21498 272662 21734
rect 272746 21498 272982 21734
rect 272426 -5382 272662 -5146
rect 272746 -5382 272982 -5146
rect 272426 -5702 272662 -5466
rect 272746 -5702 272982 -5466
rect 276146 710362 276382 710598
rect 276466 710362 276702 710598
rect 276146 710042 276382 710278
rect 276466 710042 276702 710278
rect 276146 673538 276382 673774
rect 276466 673538 276702 673774
rect 276146 673218 276382 673454
rect 276466 673218 276702 673454
rect 276146 637538 276382 637774
rect 276466 637538 276702 637774
rect 276146 637218 276382 637454
rect 276466 637218 276702 637454
rect 276146 601538 276382 601774
rect 276466 601538 276702 601774
rect 276146 601218 276382 601454
rect 276466 601218 276702 601454
rect 276146 565538 276382 565774
rect 276466 565538 276702 565774
rect 276146 565218 276382 565454
rect 276466 565218 276702 565454
rect 276146 529538 276382 529774
rect 276466 529538 276702 529774
rect 276146 529218 276382 529454
rect 276466 529218 276702 529454
rect 276146 493538 276382 493774
rect 276466 493538 276702 493774
rect 276146 493218 276382 493454
rect 276466 493218 276702 493454
rect 276146 457538 276382 457774
rect 276466 457538 276702 457774
rect 276146 457218 276382 457454
rect 276466 457218 276702 457454
rect 276146 421538 276382 421774
rect 276466 421538 276702 421774
rect 276146 421218 276382 421454
rect 276466 421218 276702 421454
rect 276146 385538 276382 385774
rect 276466 385538 276702 385774
rect 276146 385218 276382 385454
rect 276466 385218 276702 385454
rect 276146 349538 276382 349774
rect 276466 349538 276702 349774
rect 276146 349218 276382 349454
rect 276466 349218 276702 349454
rect 276146 313538 276382 313774
rect 276466 313538 276702 313774
rect 276146 313218 276382 313454
rect 276466 313218 276702 313454
rect 276146 277538 276382 277774
rect 276466 277538 276702 277774
rect 276146 277218 276382 277454
rect 276466 277218 276702 277454
rect 276146 241538 276382 241774
rect 276466 241538 276702 241774
rect 276146 241218 276382 241454
rect 276466 241218 276702 241454
rect 276146 205538 276382 205774
rect 276466 205538 276702 205774
rect 276146 205218 276382 205454
rect 276466 205218 276702 205454
rect 276146 169538 276382 169774
rect 276466 169538 276702 169774
rect 276146 169218 276382 169454
rect 276466 169218 276702 169454
rect 276146 133538 276382 133774
rect 276466 133538 276702 133774
rect 276146 133218 276382 133454
rect 276466 133218 276702 133454
rect 276146 97538 276382 97774
rect 276466 97538 276702 97774
rect 276146 97218 276382 97454
rect 276466 97218 276702 97454
rect 276146 61538 276382 61774
rect 276466 61538 276702 61774
rect 276146 61218 276382 61454
rect 276466 61218 276702 61454
rect 276146 25538 276382 25774
rect 276466 25538 276702 25774
rect 276146 25218 276382 25454
rect 276466 25218 276702 25454
rect 276146 -6342 276382 -6106
rect 276466 -6342 276702 -6106
rect 276146 -6662 276382 -6426
rect 276466 -6662 276702 -6426
rect 279866 711322 280102 711558
rect 280186 711322 280422 711558
rect 279866 711002 280102 711238
rect 280186 711002 280422 711238
rect 279866 677258 280102 677494
rect 280186 677258 280422 677494
rect 279866 676938 280102 677174
rect 280186 676938 280422 677174
rect 279866 641258 280102 641494
rect 280186 641258 280422 641494
rect 279866 640938 280102 641174
rect 280186 640938 280422 641174
rect 279866 605258 280102 605494
rect 280186 605258 280422 605494
rect 279866 604938 280102 605174
rect 280186 604938 280422 605174
rect 279866 569258 280102 569494
rect 280186 569258 280422 569494
rect 279866 568938 280102 569174
rect 280186 568938 280422 569174
rect 279866 533258 280102 533494
rect 280186 533258 280422 533494
rect 279866 532938 280102 533174
rect 280186 532938 280422 533174
rect 279866 497258 280102 497494
rect 280186 497258 280422 497494
rect 279866 496938 280102 497174
rect 280186 496938 280422 497174
rect 279866 461258 280102 461494
rect 280186 461258 280422 461494
rect 279866 460938 280102 461174
rect 280186 460938 280422 461174
rect 279866 425258 280102 425494
rect 280186 425258 280422 425494
rect 279866 424938 280102 425174
rect 280186 424938 280422 425174
rect 279866 389258 280102 389494
rect 280186 389258 280422 389494
rect 279866 388938 280102 389174
rect 280186 388938 280422 389174
rect 279866 353258 280102 353494
rect 280186 353258 280422 353494
rect 279866 352938 280102 353174
rect 280186 352938 280422 353174
rect 279866 317258 280102 317494
rect 280186 317258 280422 317494
rect 279866 316938 280102 317174
rect 280186 316938 280422 317174
rect 279866 281258 280102 281494
rect 280186 281258 280422 281494
rect 279866 280938 280102 281174
rect 280186 280938 280422 281174
rect 279866 245258 280102 245494
rect 280186 245258 280422 245494
rect 279866 244938 280102 245174
rect 280186 244938 280422 245174
rect 279866 209258 280102 209494
rect 280186 209258 280422 209494
rect 279866 208938 280102 209174
rect 280186 208938 280422 209174
rect 279866 173258 280102 173494
rect 280186 173258 280422 173494
rect 279866 172938 280102 173174
rect 280186 172938 280422 173174
rect 279866 137258 280102 137494
rect 280186 137258 280422 137494
rect 279866 136938 280102 137174
rect 280186 136938 280422 137174
rect 279866 101258 280102 101494
rect 280186 101258 280422 101494
rect 279866 100938 280102 101174
rect 280186 100938 280422 101174
rect 279866 65258 280102 65494
rect 280186 65258 280422 65494
rect 279866 64938 280102 65174
rect 280186 64938 280422 65174
rect 279866 29258 280102 29494
rect 280186 29258 280422 29494
rect 279866 28938 280102 29174
rect 280186 28938 280422 29174
rect 279866 -7302 280102 -7066
rect 280186 -7302 280422 -7066
rect 279866 -7622 280102 -7386
rect 280186 -7622 280422 -7386
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 705562 293782 705798
rect 293866 705562 294102 705798
rect 293546 705242 293782 705478
rect 293866 705242 294102 705478
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -1542 293782 -1306
rect 293866 -1542 294102 -1306
rect 293546 -1862 293782 -1626
rect 293866 -1862 294102 -1626
rect 297266 706522 297502 706758
rect 297586 706522 297822 706758
rect 297266 706202 297502 706438
rect 297586 706202 297822 706438
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -2502 297502 -2266
rect 297586 -2502 297822 -2266
rect 297266 -2822 297502 -2586
rect 297586 -2822 297822 -2586
rect 300986 707482 301222 707718
rect 301306 707482 301542 707718
rect 300986 707162 301222 707398
rect 301306 707162 301542 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 300986 -3462 301222 -3226
rect 301306 -3462 301542 -3226
rect 300986 -3782 301222 -3546
rect 301306 -3782 301542 -3546
rect 304706 708442 304942 708678
rect 305026 708442 305262 708678
rect 304706 708122 304942 708358
rect 305026 708122 305262 708358
rect 304706 666098 304942 666334
rect 305026 666098 305262 666334
rect 304706 665778 304942 666014
rect 305026 665778 305262 666014
rect 304706 630098 304942 630334
rect 305026 630098 305262 630334
rect 304706 629778 304942 630014
rect 305026 629778 305262 630014
rect 304706 594098 304942 594334
rect 305026 594098 305262 594334
rect 304706 593778 304942 594014
rect 305026 593778 305262 594014
rect 304706 558098 304942 558334
rect 305026 558098 305262 558334
rect 304706 557778 304942 558014
rect 305026 557778 305262 558014
rect 304706 522098 304942 522334
rect 305026 522098 305262 522334
rect 304706 521778 304942 522014
rect 305026 521778 305262 522014
rect 304706 486098 304942 486334
rect 305026 486098 305262 486334
rect 304706 485778 304942 486014
rect 305026 485778 305262 486014
rect 304706 450098 304942 450334
rect 305026 450098 305262 450334
rect 304706 449778 304942 450014
rect 305026 449778 305262 450014
rect 304706 414098 304942 414334
rect 305026 414098 305262 414334
rect 304706 413778 304942 414014
rect 305026 413778 305262 414014
rect 304706 378098 304942 378334
rect 305026 378098 305262 378334
rect 304706 377778 304942 378014
rect 305026 377778 305262 378014
rect 304706 342098 304942 342334
rect 305026 342098 305262 342334
rect 304706 341778 304942 342014
rect 305026 341778 305262 342014
rect 304706 306098 304942 306334
rect 305026 306098 305262 306334
rect 304706 305778 304942 306014
rect 305026 305778 305262 306014
rect 304706 270098 304942 270334
rect 305026 270098 305262 270334
rect 304706 269778 304942 270014
rect 305026 269778 305262 270014
rect 304706 234098 304942 234334
rect 305026 234098 305262 234334
rect 304706 233778 304942 234014
rect 305026 233778 305262 234014
rect 304706 198098 304942 198334
rect 305026 198098 305262 198334
rect 304706 197778 304942 198014
rect 305026 197778 305262 198014
rect 304706 162098 304942 162334
rect 305026 162098 305262 162334
rect 304706 161778 304942 162014
rect 305026 161778 305262 162014
rect 304706 126098 304942 126334
rect 305026 126098 305262 126334
rect 304706 125778 304942 126014
rect 305026 125778 305262 126014
rect 304706 90098 304942 90334
rect 305026 90098 305262 90334
rect 304706 89778 304942 90014
rect 305026 89778 305262 90014
rect 304706 54098 304942 54334
rect 305026 54098 305262 54334
rect 304706 53778 304942 54014
rect 305026 53778 305262 54014
rect 304706 18098 304942 18334
rect 305026 18098 305262 18334
rect 304706 17778 304942 18014
rect 305026 17778 305262 18014
rect 304706 -4422 304942 -4186
rect 305026 -4422 305262 -4186
rect 304706 -4742 304942 -4506
rect 305026 -4742 305262 -4506
rect 308426 709402 308662 709638
rect 308746 709402 308982 709638
rect 308426 709082 308662 709318
rect 308746 709082 308982 709318
rect 308426 669818 308662 670054
rect 308746 669818 308982 670054
rect 308426 669498 308662 669734
rect 308746 669498 308982 669734
rect 308426 633818 308662 634054
rect 308746 633818 308982 634054
rect 308426 633498 308662 633734
rect 308746 633498 308982 633734
rect 308426 597818 308662 598054
rect 308746 597818 308982 598054
rect 308426 597498 308662 597734
rect 308746 597498 308982 597734
rect 308426 561818 308662 562054
rect 308746 561818 308982 562054
rect 308426 561498 308662 561734
rect 308746 561498 308982 561734
rect 308426 525818 308662 526054
rect 308746 525818 308982 526054
rect 308426 525498 308662 525734
rect 308746 525498 308982 525734
rect 308426 489818 308662 490054
rect 308746 489818 308982 490054
rect 308426 489498 308662 489734
rect 308746 489498 308982 489734
rect 308426 453818 308662 454054
rect 308746 453818 308982 454054
rect 308426 453498 308662 453734
rect 308746 453498 308982 453734
rect 308426 417818 308662 418054
rect 308746 417818 308982 418054
rect 308426 417498 308662 417734
rect 308746 417498 308982 417734
rect 308426 381818 308662 382054
rect 308746 381818 308982 382054
rect 308426 381498 308662 381734
rect 308746 381498 308982 381734
rect 308426 345818 308662 346054
rect 308746 345818 308982 346054
rect 308426 345498 308662 345734
rect 308746 345498 308982 345734
rect 308426 309818 308662 310054
rect 308746 309818 308982 310054
rect 308426 309498 308662 309734
rect 308746 309498 308982 309734
rect 308426 273818 308662 274054
rect 308746 273818 308982 274054
rect 308426 273498 308662 273734
rect 308746 273498 308982 273734
rect 308426 237818 308662 238054
rect 308746 237818 308982 238054
rect 308426 237498 308662 237734
rect 308746 237498 308982 237734
rect 308426 201818 308662 202054
rect 308746 201818 308982 202054
rect 308426 201498 308662 201734
rect 308746 201498 308982 201734
rect 308426 165818 308662 166054
rect 308746 165818 308982 166054
rect 308426 165498 308662 165734
rect 308746 165498 308982 165734
rect 308426 129818 308662 130054
rect 308746 129818 308982 130054
rect 308426 129498 308662 129734
rect 308746 129498 308982 129734
rect 308426 93818 308662 94054
rect 308746 93818 308982 94054
rect 308426 93498 308662 93734
rect 308746 93498 308982 93734
rect 308426 57818 308662 58054
rect 308746 57818 308982 58054
rect 308426 57498 308662 57734
rect 308746 57498 308982 57734
rect 308426 21818 308662 22054
rect 308746 21818 308982 22054
rect 308426 21498 308662 21734
rect 308746 21498 308982 21734
rect 308426 -5382 308662 -5146
rect 308746 -5382 308982 -5146
rect 308426 -5702 308662 -5466
rect 308746 -5702 308982 -5466
rect 312146 710362 312382 710598
rect 312466 710362 312702 710598
rect 312146 710042 312382 710278
rect 312466 710042 312702 710278
rect 312146 673538 312382 673774
rect 312466 673538 312702 673774
rect 312146 673218 312382 673454
rect 312466 673218 312702 673454
rect 312146 637538 312382 637774
rect 312466 637538 312702 637774
rect 312146 637218 312382 637454
rect 312466 637218 312702 637454
rect 312146 601538 312382 601774
rect 312466 601538 312702 601774
rect 312146 601218 312382 601454
rect 312466 601218 312702 601454
rect 312146 565538 312382 565774
rect 312466 565538 312702 565774
rect 312146 565218 312382 565454
rect 312466 565218 312702 565454
rect 312146 529538 312382 529774
rect 312466 529538 312702 529774
rect 312146 529218 312382 529454
rect 312466 529218 312702 529454
rect 312146 493538 312382 493774
rect 312466 493538 312702 493774
rect 312146 493218 312382 493454
rect 312466 493218 312702 493454
rect 312146 457538 312382 457774
rect 312466 457538 312702 457774
rect 312146 457218 312382 457454
rect 312466 457218 312702 457454
rect 312146 421538 312382 421774
rect 312466 421538 312702 421774
rect 312146 421218 312382 421454
rect 312466 421218 312702 421454
rect 312146 385538 312382 385774
rect 312466 385538 312702 385774
rect 312146 385218 312382 385454
rect 312466 385218 312702 385454
rect 312146 349538 312382 349774
rect 312466 349538 312702 349774
rect 312146 349218 312382 349454
rect 312466 349218 312702 349454
rect 312146 313538 312382 313774
rect 312466 313538 312702 313774
rect 312146 313218 312382 313454
rect 312466 313218 312702 313454
rect 312146 277538 312382 277774
rect 312466 277538 312702 277774
rect 312146 277218 312382 277454
rect 312466 277218 312702 277454
rect 312146 241538 312382 241774
rect 312466 241538 312702 241774
rect 312146 241218 312382 241454
rect 312466 241218 312702 241454
rect 312146 205538 312382 205774
rect 312466 205538 312702 205774
rect 312146 205218 312382 205454
rect 312466 205218 312702 205454
rect 312146 169538 312382 169774
rect 312466 169538 312702 169774
rect 312146 169218 312382 169454
rect 312466 169218 312702 169454
rect 312146 133538 312382 133774
rect 312466 133538 312702 133774
rect 312146 133218 312382 133454
rect 312466 133218 312702 133454
rect 312146 97538 312382 97774
rect 312466 97538 312702 97774
rect 312146 97218 312382 97454
rect 312466 97218 312702 97454
rect 312146 61538 312382 61774
rect 312466 61538 312702 61774
rect 312146 61218 312382 61454
rect 312466 61218 312702 61454
rect 312146 25538 312382 25774
rect 312466 25538 312702 25774
rect 312146 25218 312382 25454
rect 312466 25218 312702 25454
rect 312146 -6342 312382 -6106
rect 312466 -6342 312702 -6106
rect 312146 -6662 312382 -6426
rect 312466 -6662 312702 -6426
rect 315866 711322 316102 711558
rect 316186 711322 316422 711558
rect 315866 711002 316102 711238
rect 316186 711002 316422 711238
rect 315866 677258 316102 677494
rect 316186 677258 316422 677494
rect 315866 676938 316102 677174
rect 316186 676938 316422 677174
rect 315866 641258 316102 641494
rect 316186 641258 316422 641494
rect 315866 640938 316102 641174
rect 316186 640938 316422 641174
rect 315866 605258 316102 605494
rect 316186 605258 316422 605494
rect 315866 604938 316102 605174
rect 316186 604938 316422 605174
rect 315866 569258 316102 569494
rect 316186 569258 316422 569494
rect 315866 568938 316102 569174
rect 316186 568938 316422 569174
rect 315866 533258 316102 533494
rect 316186 533258 316422 533494
rect 315866 532938 316102 533174
rect 316186 532938 316422 533174
rect 315866 497258 316102 497494
rect 316186 497258 316422 497494
rect 315866 496938 316102 497174
rect 316186 496938 316422 497174
rect 315866 461258 316102 461494
rect 316186 461258 316422 461494
rect 315866 460938 316102 461174
rect 316186 460938 316422 461174
rect 315866 425258 316102 425494
rect 316186 425258 316422 425494
rect 315866 424938 316102 425174
rect 316186 424938 316422 425174
rect 315866 389258 316102 389494
rect 316186 389258 316422 389494
rect 315866 388938 316102 389174
rect 316186 388938 316422 389174
rect 315866 353258 316102 353494
rect 316186 353258 316422 353494
rect 315866 352938 316102 353174
rect 316186 352938 316422 353174
rect 315866 317258 316102 317494
rect 316186 317258 316422 317494
rect 315866 316938 316102 317174
rect 316186 316938 316422 317174
rect 315866 281258 316102 281494
rect 316186 281258 316422 281494
rect 315866 280938 316102 281174
rect 316186 280938 316422 281174
rect 315866 245258 316102 245494
rect 316186 245258 316422 245494
rect 315866 244938 316102 245174
rect 316186 244938 316422 245174
rect 315866 209258 316102 209494
rect 316186 209258 316422 209494
rect 315866 208938 316102 209174
rect 316186 208938 316422 209174
rect 315866 173258 316102 173494
rect 316186 173258 316422 173494
rect 315866 172938 316102 173174
rect 316186 172938 316422 173174
rect 315866 137258 316102 137494
rect 316186 137258 316422 137494
rect 315866 136938 316102 137174
rect 316186 136938 316422 137174
rect 315866 101258 316102 101494
rect 316186 101258 316422 101494
rect 315866 100938 316102 101174
rect 316186 100938 316422 101174
rect 315866 65258 316102 65494
rect 316186 65258 316422 65494
rect 315866 64938 316102 65174
rect 316186 64938 316422 65174
rect 315866 29258 316102 29494
rect 316186 29258 316422 29494
rect 315866 28938 316102 29174
rect 316186 28938 316422 29174
rect 315866 -7302 316102 -7066
rect 316186 -7302 316422 -7066
rect 315866 -7622 316102 -7386
rect 316186 -7622 316422 -7386
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 705562 329782 705798
rect 329866 705562 330102 705798
rect 329546 705242 329782 705478
rect 329866 705242 330102 705478
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -1542 329782 -1306
rect 329866 -1542 330102 -1306
rect 329546 -1862 329782 -1626
rect 329866 -1862 330102 -1626
rect 333266 706522 333502 706758
rect 333586 706522 333822 706758
rect 333266 706202 333502 706438
rect 333586 706202 333822 706438
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -2502 333502 -2266
rect 333586 -2502 333822 -2266
rect 333266 -2822 333502 -2586
rect 333586 -2822 333822 -2586
rect 336986 707482 337222 707718
rect 337306 707482 337542 707718
rect 336986 707162 337222 707398
rect 337306 707162 337542 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 336986 -3462 337222 -3226
rect 337306 -3462 337542 -3226
rect 336986 -3782 337222 -3546
rect 337306 -3782 337542 -3546
rect 340706 708442 340942 708678
rect 341026 708442 341262 708678
rect 340706 708122 340942 708358
rect 341026 708122 341262 708358
rect 340706 666098 340942 666334
rect 341026 666098 341262 666334
rect 340706 665778 340942 666014
rect 341026 665778 341262 666014
rect 340706 630098 340942 630334
rect 341026 630098 341262 630334
rect 340706 629778 340942 630014
rect 341026 629778 341262 630014
rect 340706 594098 340942 594334
rect 341026 594098 341262 594334
rect 340706 593778 340942 594014
rect 341026 593778 341262 594014
rect 340706 558098 340942 558334
rect 341026 558098 341262 558334
rect 340706 557778 340942 558014
rect 341026 557778 341262 558014
rect 340706 522098 340942 522334
rect 341026 522098 341262 522334
rect 340706 521778 340942 522014
rect 341026 521778 341262 522014
rect 340706 486098 340942 486334
rect 341026 486098 341262 486334
rect 340706 485778 340942 486014
rect 341026 485778 341262 486014
rect 340706 450098 340942 450334
rect 341026 450098 341262 450334
rect 340706 449778 340942 450014
rect 341026 449778 341262 450014
rect 340706 414098 340942 414334
rect 341026 414098 341262 414334
rect 340706 413778 340942 414014
rect 341026 413778 341262 414014
rect 340706 378098 340942 378334
rect 341026 378098 341262 378334
rect 340706 377778 340942 378014
rect 341026 377778 341262 378014
rect 340706 342098 340942 342334
rect 341026 342098 341262 342334
rect 340706 341778 340942 342014
rect 341026 341778 341262 342014
rect 340706 306098 340942 306334
rect 341026 306098 341262 306334
rect 340706 305778 340942 306014
rect 341026 305778 341262 306014
rect 340706 270098 340942 270334
rect 341026 270098 341262 270334
rect 340706 269778 340942 270014
rect 341026 269778 341262 270014
rect 340706 234098 340942 234334
rect 341026 234098 341262 234334
rect 340706 233778 340942 234014
rect 341026 233778 341262 234014
rect 340706 198098 340942 198334
rect 341026 198098 341262 198334
rect 340706 197778 340942 198014
rect 341026 197778 341262 198014
rect 340706 162098 340942 162334
rect 341026 162098 341262 162334
rect 340706 161778 340942 162014
rect 341026 161778 341262 162014
rect 340706 126098 340942 126334
rect 341026 126098 341262 126334
rect 340706 125778 340942 126014
rect 341026 125778 341262 126014
rect 340706 90098 340942 90334
rect 341026 90098 341262 90334
rect 340706 89778 340942 90014
rect 341026 89778 341262 90014
rect 340706 54098 340942 54334
rect 341026 54098 341262 54334
rect 340706 53778 340942 54014
rect 341026 53778 341262 54014
rect 340706 18098 340942 18334
rect 341026 18098 341262 18334
rect 340706 17778 340942 18014
rect 341026 17778 341262 18014
rect 340706 -4422 340942 -4186
rect 341026 -4422 341262 -4186
rect 340706 -4742 340942 -4506
rect 341026 -4742 341262 -4506
rect 344426 709402 344662 709638
rect 344746 709402 344982 709638
rect 344426 709082 344662 709318
rect 344746 709082 344982 709318
rect 344426 669818 344662 670054
rect 344746 669818 344982 670054
rect 344426 669498 344662 669734
rect 344746 669498 344982 669734
rect 344426 633818 344662 634054
rect 344746 633818 344982 634054
rect 344426 633498 344662 633734
rect 344746 633498 344982 633734
rect 344426 597818 344662 598054
rect 344746 597818 344982 598054
rect 344426 597498 344662 597734
rect 344746 597498 344982 597734
rect 344426 561818 344662 562054
rect 344746 561818 344982 562054
rect 344426 561498 344662 561734
rect 344746 561498 344982 561734
rect 344426 525818 344662 526054
rect 344746 525818 344982 526054
rect 344426 525498 344662 525734
rect 344746 525498 344982 525734
rect 344426 489818 344662 490054
rect 344746 489818 344982 490054
rect 344426 489498 344662 489734
rect 344746 489498 344982 489734
rect 344426 453818 344662 454054
rect 344746 453818 344982 454054
rect 344426 453498 344662 453734
rect 344746 453498 344982 453734
rect 344426 417818 344662 418054
rect 344746 417818 344982 418054
rect 344426 417498 344662 417734
rect 344746 417498 344982 417734
rect 344426 381818 344662 382054
rect 344746 381818 344982 382054
rect 344426 381498 344662 381734
rect 344746 381498 344982 381734
rect 344426 345818 344662 346054
rect 344746 345818 344982 346054
rect 344426 345498 344662 345734
rect 344746 345498 344982 345734
rect 344426 309818 344662 310054
rect 344746 309818 344982 310054
rect 344426 309498 344662 309734
rect 344746 309498 344982 309734
rect 344426 273818 344662 274054
rect 344746 273818 344982 274054
rect 344426 273498 344662 273734
rect 344746 273498 344982 273734
rect 344426 237818 344662 238054
rect 344746 237818 344982 238054
rect 344426 237498 344662 237734
rect 344746 237498 344982 237734
rect 344426 201818 344662 202054
rect 344746 201818 344982 202054
rect 344426 201498 344662 201734
rect 344746 201498 344982 201734
rect 344426 165818 344662 166054
rect 344746 165818 344982 166054
rect 344426 165498 344662 165734
rect 344746 165498 344982 165734
rect 344426 129818 344662 130054
rect 344746 129818 344982 130054
rect 344426 129498 344662 129734
rect 344746 129498 344982 129734
rect 344426 93818 344662 94054
rect 344746 93818 344982 94054
rect 344426 93498 344662 93734
rect 344746 93498 344982 93734
rect 344426 57818 344662 58054
rect 344746 57818 344982 58054
rect 344426 57498 344662 57734
rect 344746 57498 344982 57734
rect 344426 21818 344662 22054
rect 344746 21818 344982 22054
rect 344426 21498 344662 21734
rect 344746 21498 344982 21734
rect 344426 -5382 344662 -5146
rect 344746 -5382 344982 -5146
rect 344426 -5702 344662 -5466
rect 344746 -5702 344982 -5466
rect 348146 710362 348382 710598
rect 348466 710362 348702 710598
rect 348146 710042 348382 710278
rect 348466 710042 348702 710278
rect 348146 673538 348382 673774
rect 348466 673538 348702 673774
rect 348146 673218 348382 673454
rect 348466 673218 348702 673454
rect 348146 637538 348382 637774
rect 348466 637538 348702 637774
rect 348146 637218 348382 637454
rect 348466 637218 348702 637454
rect 348146 601538 348382 601774
rect 348466 601538 348702 601774
rect 348146 601218 348382 601454
rect 348466 601218 348702 601454
rect 348146 565538 348382 565774
rect 348466 565538 348702 565774
rect 348146 565218 348382 565454
rect 348466 565218 348702 565454
rect 348146 529538 348382 529774
rect 348466 529538 348702 529774
rect 348146 529218 348382 529454
rect 348466 529218 348702 529454
rect 348146 493538 348382 493774
rect 348466 493538 348702 493774
rect 348146 493218 348382 493454
rect 348466 493218 348702 493454
rect 348146 457538 348382 457774
rect 348466 457538 348702 457774
rect 348146 457218 348382 457454
rect 348466 457218 348702 457454
rect 348146 421538 348382 421774
rect 348466 421538 348702 421774
rect 348146 421218 348382 421454
rect 348466 421218 348702 421454
rect 348146 385538 348382 385774
rect 348466 385538 348702 385774
rect 348146 385218 348382 385454
rect 348466 385218 348702 385454
rect 348146 349538 348382 349774
rect 348466 349538 348702 349774
rect 348146 349218 348382 349454
rect 348466 349218 348702 349454
rect 348146 313538 348382 313774
rect 348466 313538 348702 313774
rect 348146 313218 348382 313454
rect 348466 313218 348702 313454
rect 348146 277538 348382 277774
rect 348466 277538 348702 277774
rect 348146 277218 348382 277454
rect 348466 277218 348702 277454
rect 348146 241538 348382 241774
rect 348466 241538 348702 241774
rect 348146 241218 348382 241454
rect 348466 241218 348702 241454
rect 348146 205538 348382 205774
rect 348466 205538 348702 205774
rect 348146 205218 348382 205454
rect 348466 205218 348702 205454
rect 348146 169538 348382 169774
rect 348466 169538 348702 169774
rect 348146 169218 348382 169454
rect 348466 169218 348702 169454
rect 348146 133538 348382 133774
rect 348466 133538 348702 133774
rect 348146 133218 348382 133454
rect 348466 133218 348702 133454
rect 348146 97538 348382 97774
rect 348466 97538 348702 97774
rect 348146 97218 348382 97454
rect 348466 97218 348702 97454
rect 348146 61538 348382 61774
rect 348466 61538 348702 61774
rect 348146 61218 348382 61454
rect 348466 61218 348702 61454
rect 348146 25538 348382 25774
rect 348466 25538 348702 25774
rect 348146 25218 348382 25454
rect 348466 25218 348702 25454
rect 348146 -6342 348382 -6106
rect 348466 -6342 348702 -6106
rect 348146 -6662 348382 -6426
rect 348466 -6662 348702 -6426
rect 351866 711322 352102 711558
rect 352186 711322 352422 711558
rect 351866 711002 352102 711238
rect 352186 711002 352422 711238
rect 351866 677258 352102 677494
rect 352186 677258 352422 677494
rect 351866 676938 352102 677174
rect 352186 676938 352422 677174
rect 351866 641258 352102 641494
rect 352186 641258 352422 641494
rect 351866 640938 352102 641174
rect 352186 640938 352422 641174
rect 351866 605258 352102 605494
rect 352186 605258 352422 605494
rect 351866 604938 352102 605174
rect 352186 604938 352422 605174
rect 351866 569258 352102 569494
rect 352186 569258 352422 569494
rect 351866 568938 352102 569174
rect 352186 568938 352422 569174
rect 351866 533258 352102 533494
rect 352186 533258 352422 533494
rect 351866 532938 352102 533174
rect 352186 532938 352422 533174
rect 351866 497258 352102 497494
rect 352186 497258 352422 497494
rect 351866 496938 352102 497174
rect 352186 496938 352422 497174
rect 351866 461258 352102 461494
rect 352186 461258 352422 461494
rect 351866 460938 352102 461174
rect 352186 460938 352422 461174
rect 351866 425258 352102 425494
rect 352186 425258 352422 425494
rect 351866 424938 352102 425174
rect 352186 424938 352422 425174
rect 351866 389258 352102 389494
rect 352186 389258 352422 389494
rect 351866 388938 352102 389174
rect 352186 388938 352422 389174
rect 351866 353258 352102 353494
rect 352186 353258 352422 353494
rect 351866 352938 352102 353174
rect 352186 352938 352422 353174
rect 351866 317258 352102 317494
rect 352186 317258 352422 317494
rect 351866 316938 352102 317174
rect 352186 316938 352422 317174
rect 351866 281258 352102 281494
rect 352186 281258 352422 281494
rect 351866 280938 352102 281174
rect 352186 280938 352422 281174
rect 351866 245258 352102 245494
rect 352186 245258 352422 245494
rect 351866 244938 352102 245174
rect 352186 244938 352422 245174
rect 351866 209258 352102 209494
rect 352186 209258 352422 209494
rect 351866 208938 352102 209174
rect 352186 208938 352422 209174
rect 351866 173258 352102 173494
rect 352186 173258 352422 173494
rect 351866 172938 352102 173174
rect 352186 172938 352422 173174
rect 351866 137258 352102 137494
rect 352186 137258 352422 137494
rect 351866 136938 352102 137174
rect 352186 136938 352422 137174
rect 351866 101258 352102 101494
rect 352186 101258 352422 101494
rect 351866 100938 352102 101174
rect 352186 100938 352422 101174
rect 351866 65258 352102 65494
rect 352186 65258 352422 65494
rect 351866 64938 352102 65174
rect 352186 64938 352422 65174
rect 351866 29258 352102 29494
rect 352186 29258 352422 29494
rect 351866 28938 352102 29174
rect 352186 28938 352422 29174
rect 351866 -7302 352102 -7066
rect 352186 -7302 352422 -7066
rect 351866 -7622 352102 -7386
rect 352186 -7622 352422 -7386
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 705562 365782 705798
rect 365866 705562 366102 705798
rect 365546 705242 365782 705478
rect 365866 705242 366102 705478
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -1542 365782 -1306
rect 365866 -1542 366102 -1306
rect 365546 -1862 365782 -1626
rect 365866 -1862 366102 -1626
rect 369266 706522 369502 706758
rect 369586 706522 369822 706758
rect 369266 706202 369502 706438
rect 369586 706202 369822 706438
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -2502 369502 -2266
rect 369586 -2502 369822 -2266
rect 369266 -2822 369502 -2586
rect 369586 -2822 369822 -2586
rect 372986 707482 373222 707718
rect 373306 707482 373542 707718
rect 372986 707162 373222 707398
rect 373306 707162 373542 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 372986 -3462 373222 -3226
rect 373306 -3462 373542 -3226
rect 372986 -3782 373222 -3546
rect 373306 -3782 373542 -3546
rect 376706 708442 376942 708678
rect 377026 708442 377262 708678
rect 376706 708122 376942 708358
rect 377026 708122 377262 708358
rect 376706 666098 376942 666334
rect 377026 666098 377262 666334
rect 376706 665778 376942 666014
rect 377026 665778 377262 666014
rect 376706 630098 376942 630334
rect 377026 630098 377262 630334
rect 376706 629778 376942 630014
rect 377026 629778 377262 630014
rect 376706 594098 376942 594334
rect 377026 594098 377262 594334
rect 376706 593778 376942 594014
rect 377026 593778 377262 594014
rect 376706 558098 376942 558334
rect 377026 558098 377262 558334
rect 376706 557778 376942 558014
rect 377026 557778 377262 558014
rect 376706 522098 376942 522334
rect 377026 522098 377262 522334
rect 376706 521778 376942 522014
rect 377026 521778 377262 522014
rect 376706 486098 376942 486334
rect 377026 486098 377262 486334
rect 376706 485778 376942 486014
rect 377026 485778 377262 486014
rect 376706 450098 376942 450334
rect 377026 450098 377262 450334
rect 376706 449778 376942 450014
rect 377026 449778 377262 450014
rect 376706 414098 376942 414334
rect 377026 414098 377262 414334
rect 376706 413778 376942 414014
rect 377026 413778 377262 414014
rect 376706 378098 376942 378334
rect 377026 378098 377262 378334
rect 376706 377778 376942 378014
rect 377026 377778 377262 378014
rect 376706 342098 376942 342334
rect 377026 342098 377262 342334
rect 376706 341778 376942 342014
rect 377026 341778 377262 342014
rect 376706 306098 376942 306334
rect 377026 306098 377262 306334
rect 376706 305778 376942 306014
rect 377026 305778 377262 306014
rect 376706 270098 376942 270334
rect 377026 270098 377262 270334
rect 376706 269778 376942 270014
rect 377026 269778 377262 270014
rect 376706 234098 376942 234334
rect 377026 234098 377262 234334
rect 376706 233778 376942 234014
rect 377026 233778 377262 234014
rect 376706 198098 376942 198334
rect 377026 198098 377262 198334
rect 376706 197778 376942 198014
rect 377026 197778 377262 198014
rect 376706 162098 376942 162334
rect 377026 162098 377262 162334
rect 376706 161778 376942 162014
rect 377026 161778 377262 162014
rect 376706 126098 376942 126334
rect 377026 126098 377262 126334
rect 376706 125778 376942 126014
rect 377026 125778 377262 126014
rect 376706 90098 376942 90334
rect 377026 90098 377262 90334
rect 376706 89778 376942 90014
rect 377026 89778 377262 90014
rect 376706 54098 376942 54334
rect 377026 54098 377262 54334
rect 376706 53778 376942 54014
rect 377026 53778 377262 54014
rect 376706 18098 376942 18334
rect 377026 18098 377262 18334
rect 376706 17778 376942 18014
rect 377026 17778 377262 18014
rect 376706 -4422 376942 -4186
rect 377026 -4422 377262 -4186
rect 376706 -4742 376942 -4506
rect 377026 -4742 377262 -4506
rect 380426 709402 380662 709638
rect 380746 709402 380982 709638
rect 380426 709082 380662 709318
rect 380746 709082 380982 709318
rect 380426 669818 380662 670054
rect 380746 669818 380982 670054
rect 380426 669498 380662 669734
rect 380746 669498 380982 669734
rect 380426 633818 380662 634054
rect 380746 633818 380982 634054
rect 380426 633498 380662 633734
rect 380746 633498 380982 633734
rect 380426 597818 380662 598054
rect 380746 597818 380982 598054
rect 380426 597498 380662 597734
rect 380746 597498 380982 597734
rect 380426 561818 380662 562054
rect 380746 561818 380982 562054
rect 380426 561498 380662 561734
rect 380746 561498 380982 561734
rect 380426 525818 380662 526054
rect 380746 525818 380982 526054
rect 380426 525498 380662 525734
rect 380746 525498 380982 525734
rect 380426 489818 380662 490054
rect 380746 489818 380982 490054
rect 380426 489498 380662 489734
rect 380746 489498 380982 489734
rect 380426 453818 380662 454054
rect 380746 453818 380982 454054
rect 380426 453498 380662 453734
rect 380746 453498 380982 453734
rect 380426 417818 380662 418054
rect 380746 417818 380982 418054
rect 380426 417498 380662 417734
rect 380746 417498 380982 417734
rect 380426 381818 380662 382054
rect 380746 381818 380982 382054
rect 380426 381498 380662 381734
rect 380746 381498 380982 381734
rect 380426 345818 380662 346054
rect 380746 345818 380982 346054
rect 380426 345498 380662 345734
rect 380746 345498 380982 345734
rect 380426 309818 380662 310054
rect 380746 309818 380982 310054
rect 380426 309498 380662 309734
rect 380746 309498 380982 309734
rect 380426 273818 380662 274054
rect 380746 273818 380982 274054
rect 380426 273498 380662 273734
rect 380746 273498 380982 273734
rect 380426 237818 380662 238054
rect 380746 237818 380982 238054
rect 380426 237498 380662 237734
rect 380746 237498 380982 237734
rect 380426 201818 380662 202054
rect 380746 201818 380982 202054
rect 380426 201498 380662 201734
rect 380746 201498 380982 201734
rect 380426 165818 380662 166054
rect 380746 165818 380982 166054
rect 380426 165498 380662 165734
rect 380746 165498 380982 165734
rect 380426 129818 380662 130054
rect 380746 129818 380982 130054
rect 380426 129498 380662 129734
rect 380746 129498 380982 129734
rect 380426 93818 380662 94054
rect 380746 93818 380982 94054
rect 380426 93498 380662 93734
rect 380746 93498 380982 93734
rect 380426 57818 380662 58054
rect 380746 57818 380982 58054
rect 380426 57498 380662 57734
rect 380746 57498 380982 57734
rect 380426 21818 380662 22054
rect 380746 21818 380982 22054
rect 380426 21498 380662 21734
rect 380746 21498 380982 21734
rect 380426 -5382 380662 -5146
rect 380746 -5382 380982 -5146
rect 380426 -5702 380662 -5466
rect 380746 -5702 380982 -5466
rect 384146 710362 384382 710598
rect 384466 710362 384702 710598
rect 384146 710042 384382 710278
rect 384466 710042 384702 710278
rect 384146 673538 384382 673774
rect 384466 673538 384702 673774
rect 384146 673218 384382 673454
rect 384466 673218 384702 673454
rect 384146 637538 384382 637774
rect 384466 637538 384702 637774
rect 384146 637218 384382 637454
rect 384466 637218 384702 637454
rect 384146 601538 384382 601774
rect 384466 601538 384702 601774
rect 384146 601218 384382 601454
rect 384466 601218 384702 601454
rect 384146 565538 384382 565774
rect 384466 565538 384702 565774
rect 384146 565218 384382 565454
rect 384466 565218 384702 565454
rect 384146 529538 384382 529774
rect 384466 529538 384702 529774
rect 384146 529218 384382 529454
rect 384466 529218 384702 529454
rect 384146 493538 384382 493774
rect 384466 493538 384702 493774
rect 384146 493218 384382 493454
rect 384466 493218 384702 493454
rect 384146 457538 384382 457774
rect 384466 457538 384702 457774
rect 384146 457218 384382 457454
rect 384466 457218 384702 457454
rect 384146 421538 384382 421774
rect 384466 421538 384702 421774
rect 384146 421218 384382 421454
rect 384466 421218 384702 421454
rect 384146 385538 384382 385774
rect 384466 385538 384702 385774
rect 384146 385218 384382 385454
rect 384466 385218 384702 385454
rect 384146 349538 384382 349774
rect 384466 349538 384702 349774
rect 384146 349218 384382 349454
rect 384466 349218 384702 349454
rect 384146 313538 384382 313774
rect 384466 313538 384702 313774
rect 384146 313218 384382 313454
rect 384466 313218 384702 313454
rect 384146 277538 384382 277774
rect 384466 277538 384702 277774
rect 384146 277218 384382 277454
rect 384466 277218 384702 277454
rect 384146 241538 384382 241774
rect 384466 241538 384702 241774
rect 384146 241218 384382 241454
rect 384466 241218 384702 241454
rect 384146 205538 384382 205774
rect 384466 205538 384702 205774
rect 384146 205218 384382 205454
rect 384466 205218 384702 205454
rect 384146 169538 384382 169774
rect 384466 169538 384702 169774
rect 384146 169218 384382 169454
rect 384466 169218 384702 169454
rect 384146 133538 384382 133774
rect 384466 133538 384702 133774
rect 384146 133218 384382 133454
rect 384466 133218 384702 133454
rect 384146 97538 384382 97774
rect 384466 97538 384702 97774
rect 384146 97218 384382 97454
rect 384466 97218 384702 97454
rect 384146 61538 384382 61774
rect 384466 61538 384702 61774
rect 384146 61218 384382 61454
rect 384466 61218 384702 61454
rect 384146 25538 384382 25774
rect 384466 25538 384702 25774
rect 384146 25218 384382 25454
rect 384466 25218 384702 25454
rect 384146 -6342 384382 -6106
rect 384466 -6342 384702 -6106
rect 384146 -6662 384382 -6426
rect 384466 -6662 384702 -6426
rect 387866 711322 388102 711558
rect 388186 711322 388422 711558
rect 387866 711002 388102 711238
rect 388186 711002 388422 711238
rect 387866 677258 388102 677494
rect 388186 677258 388422 677494
rect 387866 676938 388102 677174
rect 388186 676938 388422 677174
rect 387866 641258 388102 641494
rect 388186 641258 388422 641494
rect 387866 640938 388102 641174
rect 388186 640938 388422 641174
rect 387866 605258 388102 605494
rect 388186 605258 388422 605494
rect 387866 604938 388102 605174
rect 388186 604938 388422 605174
rect 387866 569258 388102 569494
rect 388186 569258 388422 569494
rect 387866 568938 388102 569174
rect 388186 568938 388422 569174
rect 387866 533258 388102 533494
rect 388186 533258 388422 533494
rect 387866 532938 388102 533174
rect 388186 532938 388422 533174
rect 387866 497258 388102 497494
rect 388186 497258 388422 497494
rect 387866 496938 388102 497174
rect 388186 496938 388422 497174
rect 387866 461258 388102 461494
rect 388186 461258 388422 461494
rect 387866 460938 388102 461174
rect 388186 460938 388422 461174
rect 387866 425258 388102 425494
rect 388186 425258 388422 425494
rect 387866 424938 388102 425174
rect 388186 424938 388422 425174
rect 387866 389258 388102 389494
rect 388186 389258 388422 389494
rect 387866 388938 388102 389174
rect 388186 388938 388422 389174
rect 387866 353258 388102 353494
rect 388186 353258 388422 353494
rect 387866 352938 388102 353174
rect 388186 352938 388422 353174
rect 387866 317258 388102 317494
rect 388186 317258 388422 317494
rect 387866 316938 388102 317174
rect 388186 316938 388422 317174
rect 387866 281258 388102 281494
rect 388186 281258 388422 281494
rect 387866 280938 388102 281174
rect 388186 280938 388422 281174
rect 387866 245258 388102 245494
rect 388186 245258 388422 245494
rect 387866 244938 388102 245174
rect 388186 244938 388422 245174
rect 387866 209258 388102 209494
rect 388186 209258 388422 209494
rect 387866 208938 388102 209174
rect 388186 208938 388422 209174
rect 387866 173258 388102 173494
rect 388186 173258 388422 173494
rect 387866 172938 388102 173174
rect 388186 172938 388422 173174
rect 387866 137258 388102 137494
rect 388186 137258 388422 137494
rect 387866 136938 388102 137174
rect 388186 136938 388422 137174
rect 387866 101258 388102 101494
rect 388186 101258 388422 101494
rect 387866 100938 388102 101174
rect 388186 100938 388422 101174
rect 387866 65258 388102 65494
rect 388186 65258 388422 65494
rect 387866 64938 388102 65174
rect 388186 64938 388422 65174
rect 387866 29258 388102 29494
rect 388186 29258 388422 29494
rect 387866 28938 388102 29174
rect 388186 28938 388422 29174
rect 387866 -7302 388102 -7066
rect 388186 -7302 388422 -7066
rect 387866 -7622 388102 -7386
rect 388186 -7622 388422 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 705562 401782 705798
rect 401866 705562 402102 705798
rect 401546 705242 401782 705478
rect 401866 705242 402102 705478
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -1542 401782 -1306
rect 401866 -1542 402102 -1306
rect 401546 -1862 401782 -1626
rect 401866 -1862 402102 -1626
rect 405266 706522 405502 706758
rect 405586 706522 405822 706758
rect 405266 706202 405502 706438
rect 405586 706202 405822 706438
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -2502 405502 -2266
rect 405586 -2502 405822 -2266
rect 405266 -2822 405502 -2586
rect 405586 -2822 405822 -2586
rect 408986 707482 409222 707718
rect 409306 707482 409542 707718
rect 408986 707162 409222 707398
rect 409306 707162 409542 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 408986 -3462 409222 -3226
rect 409306 -3462 409542 -3226
rect 408986 -3782 409222 -3546
rect 409306 -3782 409542 -3546
rect 412706 708442 412942 708678
rect 413026 708442 413262 708678
rect 412706 708122 412942 708358
rect 413026 708122 413262 708358
rect 412706 666098 412942 666334
rect 413026 666098 413262 666334
rect 412706 665778 412942 666014
rect 413026 665778 413262 666014
rect 412706 630098 412942 630334
rect 413026 630098 413262 630334
rect 412706 629778 412942 630014
rect 413026 629778 413262 630014
rect 412706 594098 412942 594334
rect 413026 594098 413262 594334
rect 412706 593778 412942 594014
rect 413026 593778 413262 594014
rect 412706 558098 412942 558334
rect 413026 558098 413262 558334
rect 412706 557778 412942 558014
rect 413026 557778 413262 558014
rect 412706 522098 412942 522334
rect 413026 522098 413262 522334
rect 412706 521778 412942 522014
rect 413026 521778 413262 522014
rect 412706 486098 412942 486334
rect 413026 486098 413262 486334
rect 412706 485778 412942 486014
rect 413026 485778 413262 486014
rect 412706 450098 412942 450334
rect 413026 450098 413262 450334
rect 412706 449778 412942 450014
rect 413026 449778 413262 450014
rect 412706 414098 412942 414334
rect 413026 414098 413262 414334
rect 412706 413778 412942 414014
rect 413026 413778 413262 414014
rect 412706 378098 412942 378334
rect 413026 378098 413262 378334
rect 412706 377778 412942 378014
rect 413026 377778 413262 378014
rect 412706 342098 412942 342334
rect 413026 342098 413262 342334
rect 412706 341778 412942 342014
rect 413026 341778 413262 342014
rect 412706 306098 412942 306334
rect 413026 306098 413262 306334
rect 412706 305778 412942 306014
rect 413026 305778 413262 306014
rect 412706 270098 412942 270334
rect 413026 270098 413262 270334
rect 412706 269778 412942 270014
rect 413026 269778 413262 270014
rect 412706 234098 412942 234334
rect 413026 234098 413262 234334
rect 412706 233778 412942 234014
rect 413026 233778 413262 234014
rect 412706 198098 412942 198334
rect 413026 198098 413262 198334
rect 412706 197778 412942 198014
rect 413026 197778 413262 198014
rect 412706 162098 412942 162334
rect 413026 162098 413262 162334
rect 412706 161778 412942 162014
rect 413026 161778 413262 162014
rect 412706 126098 412942 126334
rect 413026 126098 413262 126334
rect 412706 125778 412942 126014
rect 413026 125778 413262 126014
rect 412706 90098 412942 90334
rect 413026 90098 413262 90334
rect 412706 89778 412942 90014
rect 413026 89778 413262 90014
rect 412706 54098 412942 54334
rect 413026 54098 413262 54334
rect 412706 53778 412942 54014
rect 413026 53778 413262 54014
rect 412706 18098 412942 18334
rect 413026 18098 413262 18334
rect 412706 17778 412942 18014
rect 413026 17778 413262 18014
rect 412706 -4422 412942 -4186
rect 413026 -4422 413262 -4186
rect 412706 -4742 412942 -4506
rect 413026 -4742 413262 -4506
rect 416426 709402 416662 709638
rect 416746 709402 416982 709638
rect 416426 709082 416662 709318
rect 416746 709082 416982 709318
rect 416426 669818 416662 670054
rect 416746 669818 416982 670054
rect 416426 669498 416662 669734
rect 416746 669498 416982 669734
rect 416426 633818 416662 634054
rect 416746 633818 416982 634054
rect 416426 633498 416662 633734
rect 416746 633498 416982 633734
rect 416426 597818 416662 598054
rect 416746 597818 416982 598054
rect 416426 597498 416662 597734
rect 416746 597498 416982 597734
rect 416426 561818 416662 562054
rect 416746 561818 416982 562054
rect 416426 561498 416662 561734
rect 416746 561498 416982 561734
rect 416426 525818 416662 526054
rect 416746 525818 416982 526054
rect 416426 525498 416662 525734
rect 416746 525498 416982 525734
rect 416426 489818 416662 490054
rect 416746 489818 416982 490054
rect 416426 489498 416662 489734
rect 416746 489498 416982 489734
rect 416426 453818 416662 454054
rect 416746 453818 416982 454054
rect 416426 453498 416662 453734
rect 416746 453498 416982 453734
rect 416426 417818 416662 418054
rect 416746 417818 416982 418054
rect 416426 417498 416662 417734
rect 416746 417498 416982 417734
rect 416426 381818 416662 382054
rect 416746 381818 416982 382054
rect 416426 381498 416662 381734
rect 416746 381498 416982 381734
rect 416426 345818 416662 346054
rect 416746 345818 416982 346054
rect 416426 345498 416662 345734
rect 416746 345498 416982 345734
rect 416426 309818 416662 310054
rect 416746 309818 416982 310054
rect 416426 309498 416662 309734
rect 416746 309498 416982 309734
rect 416426 273818 416662 274054
rect 416746 273818 416982 274054
rect 416426 273498 416662 273734
rect 416746 273498 416982 273734
rect 416426 237818 416662 238054
rect 416746 237818 416982 238054
rect 416426 237498 416662 237734
rect 416746 237498 416982 237734
rect 416426 201818 416662 202054
rect 416746 201818 416982 202054
rect 416426 201498 416662 201734
rect 416746 201498 416982 201734
rect 416426 165818 416662 166054
rect 416746 165818 416982 166054
rect 416426 165498 416662 165734
rect 416746 165498 416982 165734
rect 416426 129818 416662 130054
rect 416746 129818 416982 130054
rect 416426 129498 416662 129734
rect 416746 129498 416982 129734
rect 416426 93818 416662 94054
rect 416746 93818 416982 94054
rect 416426 93498 416662 93734
rect 416746 93498 416982 93734
rect 416426 57818 416662 58054
rect 416746 57818 416982 58054
rect 416426 57498 416662 57734
rect 416746 57498 416982 57734
rect 416426 21818 416662 22054
rect 416746 21818 416982 22054
rect 416426 21498 416662 21734
rect 416746 21498 416982 21734
rect 416426 -5382 416662 -5146
rect 416746 -5382 416982 -5146
rect 416426 -5702 416662 -5466
rect 416746 -5702 416982 -5466
rect 420146 710362 420382 710598
rect 420466 710362 420702 710598
rect 420146 710042 420382 710278
rect 420466 710042 420702 710278
rect 420146 673538 420382 673774
rect 420466 673538 420702 673774
rect 420146 673218 420382 673454
rect 420466 673218 420702 673454
rect 420146 637538 420382 637774
rect 420466 637538 420702 637774
rect 420146 637218 420382 637454
rect 420466 637218 420702 637454
rect 420146 601538 420382 601774
rect 420466 601538 420702 601774
rect 420146 601218 420382 601454
rect 420466 601218 420702 601454
rect 420146 565538 420382 565774
rect 420466 565538 420702 565774
rect 420146 565218 420382 565454
rect 420466 565218 420702 565454
rect 420146 529538 420382 529774
rect 420466 529538 420702 529774
rect 420146 529218 420382 529454
rect 420466 529218 420702 529454
rect 420146 493538 420382 493774
rect 420466 493538 420702 493774
rect 420146 493218 420382 493454
rect 420466 493218 420702 493454
rect 420146 457538 420382 457774
rect 420466 457538 420702 457774
rect 420146 457218 420382 457454
rect 420466 457218 420702 457454
rect 420146 421538 420382 421774
rect 420466 421538 420702 421774
rect 420146 421218 420382 421454
rect 420466 421218 420702 421454
rect 420146 385538 420382 385774
rect 420466 385538 420702 385774
rect 420146 385218 420382 385454
rect 420466 385218 420702 385454
rect 420146 349538 420382 349774
rect 420466 349538 420702 349774
rect 420146 349218 420382 349454
rect 420466 349218 420702 349454
rect 420146 313538 420382 313774
rect 420466 313538 420702 313774
rect 420146 313218 420382 313454
rect 420466 313218 420702 313454
rect 420146 277538 420382 277774
rect 420466 277538 420702 277774
rect 420146 277218 420382 277454
rect 420466 277218 420702 277454
rect 420146 241538 420382 241774
rect 420466 241538 420702 241774
rect 420146 241218 420382 241454
rect 420466 241218 420702 241454
rect 420146 205538 420382 205774
rect 420466 205538 420702 205774
rect 420146 205218 420382 205454
rect 420466 205218 420702 205454
rect 420146 169538 420382 169774
rect 420466 169538 420702 169774
rect 420146 169218 420382 169454
rect 420466 169218 420702 169454
rect 420146 133538 420382 133774
rect 420466 133538 420702 133774
rect 420146 133218 420382 133454
rect 420466 133218 420702 133454
rect 420146 97538 420382 97774
rect 420466 97538 420702 97774
rect 420146 97218 420382 97454
rect 420466 97218 420702 97454
rect 420146 61538 420382 61774
rect 420466 61538 420702 61774
rect 420146 61218 420382 61454
rect 420466 61218 420702 61454
rect 420146 25538 420382 25774
rect 420466 25538 420702 25774
rect 420146 25218 420382 25454
rect 420466 25218 420702 25454
rect 420146 -6342 420382 -6106
rect 420466 -6342 420702 -6106
rect 420146 -6662 420382 -6426
rect 420466 -6662 420702 -6426
rect 423866 711322 424102 711558
rect 424186 711322 424422 711558
rect 423866 711002 424102 711238
rect 424186 711002 424422 711238
rect 423866 677258 424102 677494
rect 424186 677258 424422 677494
rect 423866 676938 424102 677174
rect 424186 676938 424422 677174
rect 423866 641258 424102 641494
rect 424186 641258 424422 641494
rect 423866 640938 424102 641174
rect 424186 640938 424422 641174
rect 423866 605258 424102 605494
rect 424186 605258 424422 605494
rect 423866 604938 424102 605174
rect 424186 604938 424422 605174
rect 423866 569258 424102 569494
rect 424186 569258 424422 569494
rect 423866 568938 424102 569174
rect 424186 568938 424422 569174
rect 423866 533258 424102 533494
rect 424186 533258 424422 533494
rect 423866 532938 424102 533174
rect 424186 532938 424422 533174
rect 423866 497258 424102 497494
rect 424186 497258 424422 497494
rect 423866 496938 424102 497174
rect 424186 496938 424422 497174
rect 423866 461258 424102 461494
rect 424186 461258 424422 461494
rect 423866 460938 424102 461174
rect 424186 460938 424422 461174
rect 423866 425258 424102 425494
rect 424186 425258 424422 425494
rect 423866 424938 424102 425174
rect 424186 424938 424422 425174
rect 423866 389258 424102 389494
rect 424186 389258 424422 389494
rect 423866 388938 424102 389174
rect 424186 388938 424422 389174
rect 423866 353258 424102 353494
rect 424186 353258 424422 353494
rect 423866 352938 424102 353174
rect 424186 352938 424422 353174
rect 423866 317258 424102 317494
rect 424186 317258 424422 317494
rect 423866 316938 424102 317174
rect 424186 316938 424422 317174
rect 423866 281258 424102 281494
rect 424186 281258 424422 281494
rect 423866 280938 424102 281174
rect 424186 280938 424422 281174
rect 423866 245258 424102 245494
rect 424186 245258 424422 245494
rect 423866 244938 424102 245174
rect 424186 244938 424422 245174
rect 423866 209258 424102 209494
rect 424186 209258 424422 209494
rect 423866 208938 424102 209174
rect 424186 208938 424422 209174
rect 423866 173258 424102 173494
rect 424186 173258 424422 173494
rect 423866 172938 424102 173174
rect 424186 172938 424422 173174
rect 423866 137258 424102 137494
rect 424186 137258 424422 137494
rect 423866 136938 424102 137174
rect 424186 136938 424422 137174
rect 423866 101258 424102 101494
rect 424186 101258 424422 101494
rect 423866 100938 424102 101174
rect 424186 100938 424422 101174
rect 423866 65258 424102 65494
rect 424186 65258 424422 65494
rect 423866 64938 424102 65174
rect 424186 64938 424422 65174
rect 423866 29258 424102 29494
rect 424186 29258 424422 29494
rect 423866 28938 424102 29174
rect 424186 28938 424422 29174
rect 423866 -7302 424102 -7066
rect 424186 -7302 424422 -7066
rect 423866 -7622 424102 -7386
rect 424186 -7622 424422 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 705562 437782 705798
rect 437866 705562 438102 705798
rect 437546 705242 437782 705478
rect 437866 705242 438102 705478
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -1542 437782 -1306
rect 437866 -1542 438102 -1306
rect 437546 -1862 437782 -1626
rect 437866 -1862 438102 -1626
rect 441266 706522 441502 706758
rect 441586 706522 441822 706758
rect 441266 706202 441502 706438
rect 441586 706202 441822 706438
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -2502 441502 -2266
rect 441586 -2502 441822 -2266
rect 441266 -2822 441502 -2586
rect 441586 -2822 441822 -2586
rect 444986 707482 445222 707718
rect 445306 707482 445542 707718
rect 444986 707162 445222 707398
rect 445306 707162 445542 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 444986 -3462 445222 -3226
rect 445306 -3462 445542 -3226
rect 444986 -3782 445222 -3546
rect 445306 -3782 445542 -3546
rect 448706 708442 448942 708678
rect 449026 708442 449262 708678
rect 448706 708122 448942 708358
rect 449026 708122 449262 708358
rect 448706 666098 448942 666334
rect 449026 666098 449262 666334
rect 448706 665778 448942 666014
rect 449026 665778 449262 666014
rect 448706 630098 448942 630334
rect 449026 630098 449262 630334
rect 448706 629778 448942 630014
rect 449026 629778 449262 630014
rect 448706 594098 448942 594334
rect 449026 594098 449262 594334
rect 448706 593778 448942 594014
rect 449026 593778 449262 594014
rect 448706 558098 448942 558334
rect 449026 558098 449262 558334
rect 448706 557778 448942 558014
rect 449026 557778 449262 558014
rect 448706 522098 448942 522334
rect 449026 522098 449262 522334
rect 448706 521778 448942 522014
rect 449026 521778 449262 522014
rect 448706 486098 448942 486334
rect 449026 486098 449262 486334
rect 448706 485778 448942 486014
rect 449026 485778 449262 486014
rect 448706 450098 448942 450334
rect 449026 450098 449262 450334
rect 448706 449778 448942 450014
rect 449026 449778 449262 450014
rect 448706 414098 448942 414334
rect 449026 414098 449262 414334
rect 448706 413778 448942 414014
rect 449026 413778 449262 414014
rect 448706 378098 448942 378334
rect 449026 378098 449262 378334
rect 448706 377778 448942 378014
rect 449026 377778 449262 378014
rect 448706 342098 448942 342334
rect 449026 342098 449262 342334
rect 448706 341778 448942 342014
rect 449026 341778 449262 342014
rect 448706 306098 448942 306334
rect 449026 306098 449262 306334
rect 448706 305778 448942 306014
rect 449026 305778 449262 306014
rect 448706 270098 448942 270334
rect 449026 270098 449262 270334
rect 448706 269778 448942 270014
rect 449026 269778 449262 270014
rect 448706 234098 448942 234334
rect 449026 234098 449262 234334
rect 448706 233778 448942 234014
rect 449026 233778 449262 234014
rect 448706 198098 448942 198334
rect 449026 198098 449262 198334
rect 448706 197778 448942 198014
rect 449026 197778 449262 198014
rect 448706 162098 448942 162334
rect 449026 162098 449262 162334
rect 448706 161778 448942 162014
rect 449026 161778 449262 162014
rect 448706 126098 448942 126334
rect 449026 126098 449262 126334
rect 448706 125778 448942 126014
rect 449026 125778 449262 126014
rect 448706 90098 448942 90334
rect 449026 90098 449262 90334
rect 448706 89778 448942 90014
rect 449026 89778 449262 90014
rect 448706 54098 448942 54334
rect 449026 54098 449262 54334
rect 448706 53778 448942 54014
rect 449026 53778 449262 54014
rect 448706 18098 448942 18334
rect 449026 18098 449262 18334
rect 448706 17778 448942 18014
rect 449026 17778 449262 18014
rect 448706 -4422 448942 -4186
rect 449026 -4422 449262 -4186
rect 448706 -4742 448942 -4506
rect 449026 -4742 449262 -4506
rect 452426 709402 452662 709638
rect 452746 709402 452982 709638
rect 452426 709082 452662 709318
rect 452746 709082 452982 709318
rect 452426 669818 452662 670054
rect 452746 669818 452982 670054
rect 452426 669498 452662 669734
rect 452746 669498 452982 669734
rect 452426 633818 452662 634054
rect 452746 633818 452982 634054
rect 452426 633498 452662 633734
rect 452746 633498 452982 633734
rect 452426 597818 452662 598054
rect 452746 597818 452982 598054
rect 452426 597498 452662 597734
rect 452746 597498 452982 597734
rect 452426 561818 452662 562054
rect 452746 561818 452982 562054
rect 452426 561498 452662 561734
rect 452746 561498 452982 561734
rect 452426 525818 452662 526054
rect 452746 525818 452982 526054
rect 452426 525498 452662 525734
rect 452746 525498 452982 525734
rect 452426 489818 452662 490054
rect 452746 489818 452982 490054
rect 452426 489498 452662 489734
rect 452746 489498 452982 489734
rect 452426 453818 452662 454054
rect 452746 453818 452982 454054
rect 452426 453498 452662 453734
rect 452746 453498 452982 453734
rect 452426 417818 452662 418054
rect 452746 417818 452982 418054
rect 452426 417498 452662 417734
rect 452746 417498 452982 417734
rect 452426 381818 452662 382054
rect 452746 381818 452982 382054
rect 452426 381498 452662 381734
rect 452746 381498 452982 381734
rect 452426 345818 452662 346054
rect 452746 345818 452982 346054
rect 452426 345498 452662 345734
rect 452746 345498 452982 345734
rect 452426 309818 452662 310054
rect 452746 309818 452982 310054
rect 452426 309498 452662 309734
rect 452746 309498 452982 309734
rect 452426 273818 452662 274054
rect 452746 273818 452982 274054
rect 452426 273498 452662 273734
rect 452746 273498 452982 273734
rect 452426 237818 452662 238054
rect 452746 237818 452982 238054
rect 452426 237498 452662 237734
rect 452746 237498 452982 237734
rect 452426 201818 452662 202054
rect 452746 201818 452982 202054
rect 452426 201498 452662 201734
rect 452746 201498 452982 201734
rect 452426 165818 452662 166054
rect 452746 165818 452982 166054
rect 452426 165498 452662 165734
rect 452746 165498 452982 165734
rect 452426 129818 452662 130054
rect 452746 129818 452982 130054
rect 452426 129498 452662 129734
rect 452746 129498 452982 129734
rect 452426 93818 452662 94054
rect 452746 93818 452982 94054
rect 452426 93498 452662 93734
rect 452746 93498 452982 93734
rect 452426 57818 452662 58054
rect 452746 57818 452982 58054
rect 452426 57498 452662 57734
rect 452746 57498 452982 57734
rect 452426 21818 452662 22054
rect 452746 21818 452982 22054
rect 452426 21498 452662 21734
rect 452746 21498 452982 21734
rect 452426 -5382 452662 -5146
rect 452746 -5382 452982 -5146
rect 452426 -5702 452662 -5466
rect 452746 -5702 452982 -5466
rect 456146 710362 456382 710598
rect 456466 710362 456702 710598
rect 456146 710042 456382 710278
rect 456466 710042 456702 710278
rect 456146 673538 456382 673774
rect 456466 673538 456702 673774
rect 456146 673218 456382 673454
rect 456466 673218 456702 673454
rect 456146 637538 456382 637774
rect 456466 637538 456702 637774
rect 456146 637218 456382 637454
rect 456466 637218 456702 637454
rect 456146 601538 456382 601774
rect 456466 601538 456702 601774
rect 456146 601218 456382 601454
rect 456466 601218 456702 601454
rect 456146 565538 456382 565774
rect 456466 565538 456702 565774
rect 456146 565218 456382 565454
rect 456466 565218 456702 565454
rect 456146 529538 456382 529774
rect 456466 529538 456702 529774
rect 456146 529218 456382 529454
rect 456466 529218 456702 529454
rect 456146 493538 456382 493774
rect 456466 493538 456702 493774
rect 456146 493218 456382 493454
rect 456466 493218 456702 493454
rect 456146 457538 456382 457774
rect 456466 457538 456702 457774
rect 456146 457218 456382 457454
rect 456466 457218 456702 457454
rect 456146 421538 456382 421774
rect 456466 421538 456702 421774
rect 456146 421218 456382 421454
rect 456466 421218 456702 421454
rect 456146 385538 456382 385774
rect 456466 385538 456702 385774
rect 456146 385218 456382 385454
rect 456466 385218 456702 385454
rect 456146 349538 456382 349774
rect 456466 349538 456702 349774
rect 456146 349218 456382 349454
rect 456466 349218 456702 349454
rect 456146 313538 456382 313774
rect 456466 313538 456702 313774
rect 456146 313218 456382 313454
rect 456466 313218 456702 313454
rect 456146 277538 456382 277774
rect 456466 277538 456702 277774
rect 456146 277218 456382 277454
rect 456466 277218 456702 277454
rect 456146 241538 456382 241774
rect 456466 241538 456702 241774
rect 456146 241218 456382 241454
rect 456466 241218 456702 241454
rect 456146 205538 456382 205774
rect 456466 205538 456702 205774
rect 456146 205218 456382 205454
rect 456466 205218 456702 205454
rect 456146 169538 456382 169774
rect 456466 169538 456702 169774
rect 456146 169218 456382 169454
rect 456466 169218 456702 169454
rect 456146 133538 456382 133774
rect 456466 133538 456702 133774
rect 456146 133218 456382 133454
rect 456466 133218 456702 133454
rect 456146 97538 456382 97774
rect 456466 97538 456702 97774
rect 456146 97218 456382 97454
rect 456466 97218 456702 97454
rect 456146 61538 456382 61774
rect 456466 61538 456702 61774
rect 456146 61218 456382 61454
rect 456466 61218 456702 61454
rect 456146 25538 456382 25774
rect 456466 25538 456702 25774
rect 456146 25218 456382 25454
rect 456466 25218 456702 25454
rect 456146 -6342 456382 -6106
rect 456466 -6342 456702 -6106
rect 456146 -6662 456382 -6426
rect 456466 -6662 456702 -6426
rect 459866 711322 460102 711558
rect 460186 711322 460422 711558
rect 459866 711002 460102 711238
rect 460186 711002 460422 711238
rect 459866 677258 460102 677494
rect 460186 677258 460422 677494
rect 459866 676938 460102 677174
rect 460186 676938 460422 677174
rect 459866 641258 460102 641494
rect 460186 641258 460422 641494
rect 459866 640938 460102 641174
rect 460186 640938 460422 641174
rect 459866 605258 460102 605494
rect 460186 605258 460422 605494
rect 459866 604938 460102 605174
rect 460186 604938 460422 605174
rect 459866 569258 460102 569494
rect 460186 569258 460422 569494
rect 459866 568938 460102 569174
rect 460186 568938 460422 569174
rect 459866 533258 460102 533494
rect 460186 533258 460422 533494
rect 459866 532938 460102 533174
rect 460186 532938 460422 533174
rect 459866 497258 460102 497494
rect 460186 497258 460422 497494
rect 459866 496938 460102 497174
rect 460186 496938 460422 497174
rect 459866 461258 460102 461494
rect 460186 461258 460422 461494
rect 459866 460938 460102 461174
rect 460186 460938 460422 461174
rect 459866 425258 460102 425494
rect 460186 425258 460422 425494
rect 459866 424938 460102 425174
rect 460186 424938 460422 425174
rect 459866 389258 460102 389494
rect 460186 389258 460422 389494
rect 459866 388938 460102 389174
rect 460186 388938 460422 389174
rect 459866 353258 460102 353494
rect 460186 353258 460422 353494
rect 459866 352938 460102 353174
rect 460186 352938 460422 353174
rect 459866 317258 460102 317494
rect 460186 317258 460422 317494
rect 459866 316938 460102 317174
rect 460186 316938 460422 317174
rect 459866 281258 460102 281494
rect 460186 281258 460422 281494
rect 459866 280938 460102 281174
rect 460186 280938 460422 281174
rect 459866 245258 460102 245494
rect 460186 245258 460422 245494
rect 459866 244938 460102 245174
rect 460186 244938 460422 245174
rect 459866 209258 460102 209494
rect 460186 209258 460422 209494
rect 459866 208938 460102 209174
rect 460186 208938 460422 209174
rect 459866 173258 460102 173494
rect 460186 173258 460422 173494
rect 459866 172938 460102 173174
rect 460186 172938 460422 173174
rect 459866 137258 460102 137494
rect 460186 137258 460422 137494
rect 459866 136938 460102 137174
rect 460186 136938 460422 137174
rect 459866 101258 460102 101494
rect 460186 101258 460422 101494
rect 459866 100938 460102 101174
rect 460186 100938 460422 101174
rect 459866 65258 460102 65494
rect 460186 65258 460422 65494
rect 459866 64938 460102 65174
rect 460186 64938 460422 65174
rect 459866 29258 460102 29494
rect 460186 29258 460422 29494
rect 459866 28938 460102 29174
rect 460186 28938 460422 29174
rect 459866 -7302 460102 -7066
rect 460186 -7302 460422 -7066
rect 459866 -7622 460102 -7386
rect 460186 -7622 460422 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 705562 473782 705798
rect 473866 705562 474102 705798
rect 473546 705242 473782 705478
rect 473866 705242 474102 705478
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -1542 473782 -1306
rect 473866 -1542 474102 -1306
rect 473546 -1862 473782 -1626
rect 473866 -1862 474102 -1626
rect 477266 706522 477502 706758
rect 477586 706522 477822 706758
rect 477266 706202 477502 706438
rect 477586 706202 477822 706438
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -2502 477502 -2266
rect 477586 -2502 477822 -2266
rect 477266 -2822 477502 -2586
rect 477586 -2822 477822 -2586
rect 480986 707482 481222 707718
rect 481306 707482 481542 707718
rect 480986 707162 481222 707398
rect 481306 707162 481542 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 480986 -3462 481222 -3226
rect 481306 -3462 481542 -3226
rect 480986 -3782 481222 -3546
rect 481306 -3782 481542 -3546
rect 484706 708442 484942 708678
rect 485026 708442 485262 708678
rect 484706 708122 484942 708358
rect 485026 708122 485262 708358
rect 484706 666098 484942 666334
rect 485026 666098 485262 666334
rect 484706 665778 484942 666014
rect 485026 665778 485262 666014
rect 484706 630098 484942 630334
rect 485026 630098 485262 630334
rect 484706 629778 484942 630014
rect 485026 629778 485262 630014
rect 484706 594098 484942 594334
rect 485026 594098 485262 594334
rect 484706 593778 484942 594014
rect 485026 593778 485262 594014
rect 484706 558098 484942 558334
rect 485026 558098 485262 558334
rect 484706 557778 484942 558014
rect 485026 557778 485262 558014
rect 484706 522098 484942 522334
rect 485026 522098 485262 522334
rect 484706 521778 484942 522014
rect 485026 521778 485262 522014
rect 484706 486098 484942 486334
rect 485026 486098 485262 486334
rect 484706 485778 484942 486014
rect 485026 485778 485262 486014
rect 484706 450098 484942 450334
rect 485026 450098 485262 450334
rect 484706 449778 484942 450014
rect 485026 449778 485262 450014
rect 484706 414098 484942 414334
rect 485026 414098 485262 414334
rect 484706 413778 484942 414014
rect 485026 413778 485262 414014
rect 484706 378098 484942 378334
rect 485026 378098 485262 378334
rect 484706 377778 484942 378014
rect 485026 377778 485262 378014
rect 484706 342098 484942 342334
rect 485026 342098 485262 342334
rect 484706 341778 484942 342014
rect 485026 341778 485262 342014
rect 484706 306098 484942 306334
rect 485026 306098 485262 306334
rect 484706 305778 484942 306014
rect 485026 305778 485262 306014
rect 484706 270098 484942 270334
rect 485026 270098 485262 270334
rect 484706 269778 484942 270014
rect 485026 269778 485262 270014
rect 484706 234098 484942 234334
rect 485026 234098 485262 234334
rect 484706 233778 484942 234014
rect 485026 233778 485262 234014
rect 484706 198098 484942 198334
rect 485026 198098 485262 198334
rect 484706 197778 484942 198014
rect 485026 197778 485262 198014
rect 484706 162098 484942 162334
rect 485026 162098 485262 162334
rect 484706 161778 484942 162014
rect 485026 161778 485262 162014
rect 484706 126098 484942 126334
rect 485026 126098 485262 126334
rect 484706 125778 484942 126014
rect 485026 125778 485262 126014
rect 484706 90098 484942 90334
rect 485026 90098 485262 90334
rect 484706 89778 484942 90014
rect 485026 89778 485262 90014
rect 484706 54098 484942 54334
rect 485026 54098 485262 54334
rect 484706 53778 484942 54014
rect 485026 53778 485262 54014
rect 484706 18098 484942 18334
rect 485026 18098 485262 18334
rect 484706 17778 484942 18014
rect 485026 17778 485262 18014
rect 484706 -4422 484942 -4186
rect 485026 -4422 485262 -4186
rect 484706 -4742 484942 -4506
rect 485026 -4742 485262 -4506
rect 488426 709402 488662 709638
rect 488746 709402 488982 709638
rect 488426 709082 488662 709318
rect 488746 709082 488982 709318
rect 488426 669818 488662 670054
rect 488746 669818 488982 670054
rect 488426 669498 488662 669734
rect 488746 669498 488982 669734
rect 488426 633818 488662 634054
rect 488746 633818 488982 634054
rect 488426 633498 488662 633734
rect 488746 633498 488982 633734
rect 488426 597818 488662 598054
rect 488746 597818 488982 598054
rect 488426 597498 488662 597734
rect 488746 597498 488982 597734
rect 488426 561818 488662 562054
rect 488746 561818 488982 562054
rect 488426 561498 488662 561734
rect 488746 561498 488982 561734
rect 488426 525818 488662 526054
rect 488746 525818 488982 526054
rect 488426 525498 488662 525734
rect 488746 525498 488982 525734
rect 488426 489818 488662 490054
rect 488746 489818 488982 490054
rect 488426 489498 488662 489734
rect 488746 489498 488982 489734
rect 488426 453818 488662 454054
rect 488746 453818 488982 454054
rect 488426 453498 488662 453734
rect 488746 453498 488982 453734
rect 488426 417818 488662 418054
rect 488746 417818 488982 418054
rect 488426 417498 488662 417734
rect 488746 417498 488982 417734
rect 488426 381818 488662 382054
rect 488746 381818 488982 382054
rect 488426 381498 488662 381734
rect 488746 381498 488982 381734
rect 488426 345818 488662 346054
rect 488746 345818 488982 346054
rect 488426 345498 488662 345734
rect 488746 345498 488982 345734
rect 488426 309818 488662 310054
rect 488746 309818 488982 310054
rect 488426 309498 488662 309734
rect 488746 309498 488982 309734
rect 488426 273818 488662 274054
rect 488746 273818 488982 274054
rect 488426 273498 488662 273734
rect 488746 273498 488982 273734
rect 488426 237818 488662 238054
rect 488746 237818 488982 238054
rect 488426 237498 488662 237734
rect 488746 237498 488982 237734
rect 488426 201818 488662 202054
rect 488746 201818 488982 202054
rect 488426 201498 488662 201734
rect 488746 201498 488982 201734
rect 488426 165818 488662 166054
rect 488746 165818 488982 166054
rect 488426 165498 488662 165734
rect 488746 165498 488982 165734
rect 488426 129818 488662 130054
rect 488746 129818 488982 130054
rect 488426 129498 488662 129734
rect 488746 129498 488982 129734
rect 488426 93818 488662 94054
rect 488746 93818 488982 94054
rect 488426 93498 488662 93734
rect 488746 93498 488982 93734
rect 488426 57818 488662 58054
rect 488746 57818 488982 58054
rect 488426 57498 488662 57734
rect 488746 57498 488982 57734
rect 488426 21818 488662 22054
rect 488746 21818 488982 22054
rect 488426 21498 488662 21734
rect 488746 21498 488982 21734
rect 488426 -5382 488662 -5146
rect 488746 -5382 488982 -5146
rect 488426 -5702 488662 -5466
rect 488746 -5702 488982 -5466
rect 492146 710362 492382 710598
rect 492466 710362 492702 710598
rect 492146 710042 492382 710278
rect 492466 710042 492702 710278
rect 492146 673538 492382 673774
rect 492466 673538 492702 673774
rect 492146 673218 492382 673454
rect 492466 673218 492702 673454
rect 492146 637538 492382 637774
rect 492466 637538 492702 637774
rect 492146 637218 492382 637454
rect 492466 637218 492702 637454
rect 492146 601538 492382 601774
rect 492466 601538 492702 601774
rect 492146 601218 492382 601454
rect 492466 601218 492702 601454
rect 492146 565538 492382 565774
rect 492466 565538 492702 565774
rect 492146 565218 492382 565454
rect 492466 565218 492702 565454
rect 492146 529538 492382 529774
rect 492466 529538 492702 529774
rect 492146 529218 492382 529454
rect 492466 529218 492702 529454
rect 492146 493538 492382 493774
rect 492466 493538 492702 493774
rect 492146 493218 492382 493454
rect 492466 493218 492702 493454
rect 492146 457538 492382 457774
rect 492466 457538 492702 457774
rect 492146 457218 492382 457454
rect 492466 457218 492702 457454
rect 492146 421538 492382 421774
rect 492466 421538 492702 421774
rect 492146 421218 492382 421454
rect 492466 421218 492702 421454
rect 492146 385538 492382 385774
rect 492466 385538 492702 385774
rect 492146 385218 492382 385454
rect 492466 385218 492702 385454
rect 492146 349538 492382 349774
rect 492466 349538 492702 349774
rect 492146 349218 492382 349454
rect 492466 349218 492702 349454
rect 492146 313538 492382 313774
rect 492466 313538 492702 313774
rect 492146 313218 492382 313454
rect 492466 313218 492702 313454
rect 492146 277538 492382 277774
rect 492466 277538 492702 277774
rect 492146 277218 492382 277454
rect 492466 277218 492702 277454
rect 492146 241538 492382 241774
rect 492466 241538 492702 241774
rect 492146 241218 492382 241454
rect 492466 241218 492702 241454
rect 492146 205538 492382 205774
rect 492466 205538 492702 205774
rect 492146 205218 492382 205454
rect 492466 205218 492702 205454
rect 492146 169538 492382 169774
rect 492466 169538 492702 169774
rect 492146 169218 492382 169454
rect 492466 169218 492702 169454
rect 492146 133538 492382 133774
rect 492466 133538 492702 133774
rect 492146 133218 492382 133454
rect 492466 133218 492702 133454
rect 492146 97538 492382 97774
rect 492466 97538 492702 97774
rect 492146 97218 492382 97454
rect 492466 97218 492702 97454
rect 492146 61538 492382 61774
rect 492466 61538 492702 61774
rect 492146 61218 492382 61454
rect 492466 61218 492702 61454
rect 492146 25538 492382 25774
rect 492466 25538 492702 25774
rect 492146 25218 492382 25454
rect 492466 25218 492702 25454
rect 492146 -6342 492382 -6106
rect 492466 -6342 492702 -6106
rect 492146 -6662 492382 -6426
rect 492466 -6662 492702 -6426
rect 495866 711322 496102 711558
rect 496186 711322 496422 711558
rect 495866 711002 496102 711238
rect 496186 711002 496422 711238
rect 495866 677258 496102 677494
rect 496186 677258 496422 677494
rect 495866 676938 496102 677174
rect 496186 676938 496422 677174
rect 495866 641258 496102 641494
rect 496186 641258 496422 641494
rect 495866 640938 496102 641174
rect 496186 640938 496422 641174
rect 495866 605258 496102 605494
rect 496186 605258 496422 605494
rect 495866 604938 496102 605174
rect 496186 604938 496422 605174
rect 495866 569258 496102 569494
rect 496186 569258 496422 569494
rect 495866 568938 496102 569174
rect 496186 568938 496422 569174
rect 495866 533258 496102 533494
rect 496186 533258 496422 533494
rect 495866 532938 496102 533174
rect 496186 532938 496422 533174
rect 495866 497258 496102 497494
rect 496186 497258 496422 497494
rect 495866 496938 496102 497174
rect 496186 496938 496422 497174
rect 495866 461258 496102 461494
rect 496186 461258 496422 461494
rect 495866 460938 496102 461174
rect 496186 460938 496422 461174
rect 495866 425258 496102 425494
rect 496186 425258 496422 425494
rect 495866 424938 496102 425174
rect 496186 424938 496422 425174
rect 495866 389258 496102 389494
rect 496186 389258 496422 389494
rect 495866 388938 496102 389174
rect 496186 388938 496422 389174
rect 495866 353258 496102 353494
rect 496186 353258 496422 353494
rect 495866 352938 496102 353174
rect 496186 352938 496422 353174
rect 495866 317258 496102 317494
rect 496186 317258 496422 317494
rect 495866 316938 496102 317174
rect 496186 316938 496422 317174
rect 495866 281258 496102 281494
rect 496186 281258 496422 281494
rect 495866 280938 496102 281174
rect 496186 280938 496422 281174
rect 495866 245258 496102 245494
rect 496186 245258 496422 245494
rect 495866 244938 496102 245174
rect 496186 244938 496422 245174
rect 495866 209258 496102 209494
rect 496186 209258 496422 209494
rect 495866 208938 496102 209174
rect 496186 208938 496422 209174
rect 495866 173258 496102 173494
rect 496186 173258 496422 173494
rect 495866 172938 496102 173174
rect 496186 172938 496422 173174
rect 495866 137258 496102 137494
rect 496186 137258 496422 137494
rect 495866 136938 496102 137174
rect 496186 136938 496422 137174
rect 495866 101258 496102 101494
rect 496186 101258 496422 101494
rect 495866 100938 496102 101174
rect 496186 100938 496422 101174
rect 495866 65258 496102 65494
rect 496186 65258 496422 65494
rect 495866 64938 496102 65174
rect 496186 64938 496422 65174
rect 495866 29258 496102 29494
rect 496186 29258 496422 29494
rect 495866 28938 496102 29174
rect 496186 28938 496422 29174
rect 495866 -7302 496102 -7066
rect 496186 -7302 496422 -7066
rect 495866 -7622 496102 -7386
rect 496186 -7622 496422 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 705562 509782 705798
rect 509866 705562 510102 705798
rect 509546 705242 509782 705478
rect 509866 705242 510102 705478
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -1542 509782 -1306
rect 509866 -1542 510102 -1306
rect 509546 -1862 509782 -1626
rect 509866 -1862 510102 -1626
rect 513266 706522 513502 706758
rect 513586 706522 513822 706758
rect 513266 706202 513502 706438
rect 513586 706202 513822 706438
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -2502 513502 -2266
rect 513586 -2502 513822 -2266
rect 513266 -2822 513502 -2586
rect 513586 -2822 513822 -2586
rect 516986 707482 517222 707718
rect 517306 707482 517542 707718
rect 516986 707162 517222 707398
rect 517306 707162 517542 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 516986 -3462 517222 -3226
rect 517306 -3462 517542 -3226
rect 516986 -3782 517222 -3546
rect 517306 -3782 517542 -3546
rect 520706 708442 520942 708678
rect 521026 708442 521262 708678
rect 520706 708122 520942 708358
rect 521026 708122 521262 708358
rect 520706 666098 520942 666334
rect 521026 666098 521262 666334
rect 520706 665778 520942 666014
rect 521026 665778 521262 666014
rect 520706 630098 520942 630334
rect 521026 630098 521262 630334
rect 520706 629778 520942 630014
rect 521026 629778 521262 630014
rect 520706 594098 520942 594334
rect 521026 594098 521262 594334
rect 520706 593778 520942 594014
rect 521026 593778 521262 594014
rect 520706 558098 520942 558334
rect 521026 558098 521262 558334
rect 520706 557778 520942 558014
rect 521026 557778 521262 558014
rect 520706 522098 520942 522334
rect 521026 522098 521262 522334
rect 520706 521778 520942 522014
rect 521026 521778 521262 522014
rect 520706 486098 520942 486334
rect 521026 486098 521262 486334
rect 520706 485778 520942 486014
rect 521026 485778 521262 486014
rect 520706 450098 520942 450334
rect 521026 450098 521262 450334
rect 520706 449778 520942 450014
rect 521026 449778 521262 450014
rect 520706 414098 520942 414334
rect 521026 414098 521262 414334
rect 520706 413778 520942 414014
rect 521026 413778 521262 414014
rect 520706 378098 520942 378334
rect 521026 378098 521262 378334
rect 520706 377778 520942 378014
rect 521026 377778 521262 378014
rect 520706 342098 520942 342334
rect 521026 342098 521262 342334
rect 520706 341778 520942 342014
rect 521026 341778 521262 342014
rect 520706 306098 520942 306334
rect 521026 306098 521262 306334
rect 520706 305778 520942 306014
rect 521026 305778 521262 306014
rect 520706 270098 520942 270334
rect 521026 270098 521262 270334
rect 520706 269778 520942 270014
rect 521026 269778 521262 270014
rect 520706 234098 520942 234334
rect 521026 234098 521262 234334
rect 520706 233778 520942 234014
rect 521026 233778 521262 234014
rect 520706 198098 520942 198334
rect 521026 198098 521262 198334
rect 520706 197778 520942 198014
rect 521026 197778 521262 198014
rect 520706 162098 520942 162334
rect 521026 162098 521262 162334
rect 520706 161778 520942 162014
rect 521026 161778 521262 162014
rect 520706 126098 520942 126334
rect 521026 126098 521262 126334
rect 520706 125778 520942 126014
rect 521026 125778 521262 126014
rect 520706 90098 520942 90334
rect 521026 90098 521262 90334
rect 520706 89778 520942 90014
rect 521026 89778 521262 90014
rect 520706 54098 520942 54334
rect 521026 54098 521262 54334
rect 520706 53778 520942 54014
rect 521026 53778 521262 54014
rect 520706 18098 520942 18334
rect 521026 18098 521262 18334
rect 520706 17778 520942 18014
rect 521026 17778 521262 18014
rect 520706 -4422 520942 -4186
rect 521026 -4422 521262 -4186
rect 520706 -4742 520942 -4506
rect 521026 -4742 521262 -4506
rect 524426 709402 524662 709638
rect 524746 709402 524982 709638
rect 524426 709082 524662 709318
rect 524746 709082 524982 709318
rect 524426 669818 524662 670054
rect 524746 669818 524982 670054
rect 524426 669498 524662 669734
rect 524746 669498 524982 669734
rect 524426 633818 524662 634054
rect 524746 633818 524982 634054
rect 524426 633498 524662 633734
rect 524746 633498 524982 633734
rect 524426 597818 524662 598054
rect 524746 597818 524982 598054
rect 524426 597498 524662 597734
rect 524746 597498 524982 597734
rect 524426 561818 524662 562054
rect 524746 561818 524982 562054
rect 524426 561498 524662 561734
rect 524746 561498 524982 561734
rect 524426 525818 524662 526054
rect 524746 525818 524982 526054
rect 524426 525498 524662 525734
rect 524746 525498 524982 525734
rect 524426 489818 524662 490054
rect 524746 489818 524982 490054
rect 524426 489498 524662 489734
rect 524746 489498 524982 489734
rect 524426 453818 524662 454054
rect 524746 453818 524982 454054
rect 524426 453498 524662 453734
rect 524746 453498 524982 453734
rect 524426 417818 524662 418054
rect 524746 417818 524982 418054
rect 524426 417498 524662 417734
rect 524746 417498 524982 417734
rect 524426 381818 524662 382054
rect 524746 381818 524982 382054
rect 524426 381498 524662 381734
rect 524746 381498 524982 381734
rect 524426 345818 524662 346054
rect 524746 345818 524982 346054
rect 524426 345498 524662 345734
rect 524746 345498 524982 345734
rect 524426 309818 524662 310054
rect 524746 309818 524982 310054
rect 524426 309498 524662 309734
rect 524746 309498 524982 309734
rect 524426 273818 524662 274054
rect 524746 273818 524982 274054
rect 524426 273498 524662 273734
rect 524746 273498 524982 273734
rect 524426 237818 524662 238054
rect 524746 237818 524982 238054
rect 524426 237498 524662 237734
rect 524746 237498 524982 237734
rect 524426 201818 524662 202054
rect 524746 201818 524982 202054
rect 524426 201498 524662 201734
rect 524746 201498 524982 201734
rect 524426 165818 524662 166054
rect 524746 165818 524982 166054
rect 524426 165498 524662 165734
rect 524746 165498 524982 165734
rect 524426 129818 524662 130054
rect 524746 129818 524982 130054
rect 524426 129498 524662 129734
rect 524746 129498 524982 129734
rect 524426 93818 524662 94054
rect 524746 93818 524982 94054
rect 524426 93498 524662 93734
rect 524746 93498 524982 93734
rect 524426 57818 524662 58054
rect 524746 57818 524982 58054
rect 524426 57498 524662 57734
rect 524746 57498 524982 57734
rect 524426 21818 524662 22054
rect 524746 21818 524982 22054
rect 524426 21498 524662 21734
rect 524746 21498 524982 21734
rect 524426 -5382 524662 -5146
rect 524746 -5382 524982 -5146
rect 524426 -5702 524662 -5466
rect 524746 -5702 524982 -5466
rect 528146 710362 528382 710598
rect 528466 710362 528702 710598
rect 528146 710042 528382 710278
rect 528466 710042 528702 710278
rect 528146 673538 528382 673774
rect 528466 673538 528702 673774
rect 528146 673218 528382 673454
rect 528466 673218 528702 673454
rect 528146 637538 528382 637774
rect 528466 637538 528702 637774
rect 528146 637218 528382 637454
rect 528466 637218 528702 637454
rect 528146 601538 528382 601774
rect 528466 601538 528702 601774
rect 528146 601218 528382 601454
rect 528466 601218 528702 601454
rect 528146 565538 528382 565774
rect 528466 565538 528702 565774
rect 528146 565218 528382 565454
rect 528466 565218 528702 565454
rect 528146 529538 528382 529774
rect 528466 529538 528702 529774
rect 528146 529218 528382 529454
rect 528466 529218 528702 529454
rect 528146 493538 528382 493774
rect 528466 493538 528702 493774
rect 528146 493218 528382 493454
rect 528466 493218 528702 493454
rect 528146 457538 528382 457774
rect 528466 457538 528702 457774
rect 528146 457218 528382 457454
rect 528466 457218 528702 457454
rect 528146 421538 528382 421774
rect 528466 421538 528702 421774
rect 528146 421218 528382 421454
rect 528466 421218 528702 421454
rect 528146 385538 528382 385774
rect 528466 385538 528702 385774
rect 528146 385218 528382 385454
rect 528466 385218 528702 385454
rect 528146 349538 528382 349774
rect 528466 349538 528702 349774
rect 528146 349218 528382 349454
rect 528466 349218 528702 349454
rect 528146 313538 528382 313774
rect 528466 313538 528702 313774
rect 528146 313218 528382 313454
rect 528466 313218 528702 313454
rect 528146 277538 528382 277774
rect 528466 277538 528702 277774
rect 528146 277218 528382 277454
rect 528466 277218 528702 277454
rect 528146 241538 528382 241774
rect 528466 241538 528702 241774
rect 528146 241218 528382 241454
rect 528466 241218 528702 241454
rect 528146 205538 528382 205774
rect 528466 205538 528702 205774
rect 528146 205218 528382 205454
rect 528466 205218 528702 205454
rect 528146 169538 528382 169774
rect 528466 169538 528702 169774
rect 528146 169218 528382 169454
rect 528466 169218 528702 169454
rect 528146 133538 528382 133774
rect 528466 133538 528702 133774
rect 528146 133218 528382 133454
rect 528466 133218 528702 133454
rect 528146 97538 528382 97774
rect 528466 97538 528702 97774
rect 528146 97218 528382 97454
rect 528466 97218 528702 97454
rect 528146 61538 528382 61774
rect 528466 61538 528702 61774
rect 528146 61218 528382 61454
rect 528466 61218 528702 61454
rect 528146 25538 528382 25774
rect 528466 25538 528702 25774
rect 528146 25218 528382 25454
rect 528466 25218 528702 25454
rect 528146 -6342 528382 -6106
rect 528466 -6342 528702 -6106
rect 528146 -6662 528382 -6426
rect 528466 -6662 528702 -6426
rect 531866 711322 532102 711558
rect 532186 711322 532422 711558
rect 531866 711002 532102 711238
rect 532186 711002 532422 711238
rect 531866 677258 532102 677494
rect 532186 677258 532422 677494
rect 531866 676938 532102 677174
rect 532186 676938 532422 677174
rect 531866 641258 532102 641494
rect 532186 641258 532422 641494
rect 531866 640938 532102 641174
rect 532186 640938 532422 641174
rect 531866 605258 532102 605494
rect 532186 605258 532422 605494
rect 531866 604938 532102 605174
rect 532186 604938 532422 605174
rect 531866 569258 532102 569494
rect 532186 569258 532422 569494
rect 531866 568938 532102 569174
rect 532186 568938 532422 569174
rect 531866 533258 532102 533494
rect 532186 533258 532422 533494
rect 531866 532938 532102 533174
rect 532186 532938 532422 533174
rect 531866 497258 532102 497494
rect 532186 497258 532422 497494
rect 531866 496938 532102 497174
rect 532186 496938 532422 497174
rect 531866 461258 532102 461494
rect 532186 461258 532422 461494
rect 531866 460938 532102 461174
rect 532186 460938 532422 461174
rect 531866 425258 532102 425494
rect 532186 425258 532422 425494
rect 531866 424938 532102 425174
rect 532186 424938 532422 425174
rect 531866 389258 532102 389494
rect 532186 389258 532422 389494
rect 531866 388938 532102 389174
rect 532186 388938 532422 389174
rect 531866 353258 532102 353494
rect 532186 353258 532422 353494
rect 531866 352938 532102 353174
rect 532186 352938 532422 353174
rect 531866 317258 532102 317494
rect 532186 317258 532422 317494
rect 531866 316938 532102 317174
rect 532186 316938 532422 317174
rect 531866 281258 532102 281494
rect 532186 281258 532422 281494
rect 531866 280938 532102 281174
rect 532186 280938 532422 281174
rect 531866 245258 532102 245494
rect 532186 245258 532422 245494
rect 531866 244938 532102 245174
rect 532186 244938 532422 245174
rect 531866 209258 532102 209494
rect 532186 209258 532422 209494
rect 531866 208938 532102 209174
rect 532186 208938 532422 209174
rect 531866 173258 532102 173494
rect 532186 173258 532422 173494
rect 531866 172938 532102 173174
rect 532186 172938 532422 173174
rect 531866 137258 532102 137494
rect 532186 137258 532422 137494
rect 531866 136938 532102 137174
rect 532186 136938 532422 137174
rect 531866 101258 532102 101494
rect 532186 101258 532422 101494
rect 531866 100938 532102 101174
rect 532186 100938 532422 101174
rect 531866 65258 532102 65494
rect 532186 65258 532422 65494
rect 531866 64938 532102 65174
rect 532186 64938 532422 65174
rect 531866 29258 532102 29494
rect 532186 29258 532422 29494
rect 531866 28938 532102 29174
rect 532186 28938 532422 29174
rect 531866 -7302 532102 -7066
rect 532186 -7302 532422 -7066
rect 531866 -7622 532102 -7386
rect 532186 -7622 532422 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 705562 545782 705798
rect 545866 705562 546102 705798
rect 545546 705242 545782 705478
rect 545866 705242 546102 705478
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -1542 545782 -1306
rect 545866 -1542 546102 -1306
rect 545546 -1862 545782 -1626
rect 545866 -1862 546102 -1626
rect 549266 706522 549502 706758
rect 549586 706522 549822 706758
rect 549266 706202 549502 706438
rect 549586 706202 549822 706438
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -2502 549502 -2266
rect 549586 -2502 549822 -2266
rect 549266 -2822 549502 -2586
rect 549586 -2822 549822 -2586
rect 552986 707482 553222 707718
rect 553306 707482 553542 707718
rect 552986 707162 553222 707398
rect 553306 707162 553542 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 552986 -3462 553222 -3226
rect 553306 -3462 553542 -3226
rect 552986 -3782 553222 -3546
rect 553306 -3782 553542 -3546
rect 556706 708442 556942 708678
rect 557026 708442 557262 708678
rect 556706 708122 556942 708358
rect 557026 708122 557262 708358
rect 556706 666098 556942 666334
rect 557026 666098 557262 666334
rect 556706 665778 556942 666014
rect 557026 665778 557262 666014
rect 556706 630098 556942 630334
rect 557026 630098 557262 630334
rect 556706 629778 556942 630014
rect 557026 629778 557262 630014
rect 556706 594098 556942 594334
rect 557026 594098 557262 594334
rect 556706 593778 556942 594014
rect 557026 593778 557262 594014
rect 556706 558098 556942 558334
rect 557026 558098 557262 558334
rect 556706 557778 556942 558014
rect 557026 557778 557262 558014
rect 556706 522098 556942 522334
rect 557026 522098 557262 522334
rect 556706 521778 556942 522014
rect 557026 521778 557262 522014
rect 556706 486098 556942 486334
rect 557026 486098 557262 486334
rect 556706 485778 556942 486014
rect 557026 485778 557262 486014
rect 556706 450098 556942 450334
rect 557026 450098 557262 450334
rect 556706 449778 556942 450014
rect 557026 449778 557262 450014
rect 556706 414098 556942 414334
rect 557026 414098 557262 414334
rect 556706 413778 556942 414014
rect 557026 413778 557262 414014
rect 556706 378098 556942 378334
rect 557026 378098 557262 378334
rect 556706 377778 556942 378014
rect 557026 377778 557262 378014
rect 556706 342098 556942 342334
rect 557026 342098 557262 342334
rect 556706 341778 556942 342014
rect 557026 341778 557262 342014
rect 556706 306098 556942 306334
rect 557026 306098 557262 306334
rect 556706 305778 556942 306014
rect 557026 305778 557262 306014
rect 556706 270098 556942 270334
rect 557026 270098 557262 270334
rect 556706 269778 556942 270014
rect 557026 269778 557262 270014
rect 556706 234098 556942 234334
rect 557026 234098 557262 234334
rect 556706 233778 556942 234014
rect 557026 233778 557262 234014
rect 556706 198098 556942 198334
rect 557026 198098 557262 198334
rect 556706 197778 556942 198014
rect 557026 197778 557262 198014
rect 556706 162098 556942 162334
rect 557026 162098 557262 162334
rect 556706 161778 556942 162014
rect 557026 161778 557262 162014
rect 556706 126098 556942 126334
rect 557026 126098 557262 126334
rect 556706 125778 556942 126014
rect 557026 125778 557262 126014
rect 556706 90098 556942 90334
rect 557026 90098 557262 90334
rect 556706 89778 556942 90014
rect 557026 89778 557262 90014
rect 556706 54098 556942 54334
rect 557026 54098 557262 54334
rect 556706 53778 556942 54014
rect 557026 53778 557262 54014
rect 556706 18098 556942 18334
rect 557026 18098 557262 18334
rect 556706 17778 556942 18014
rect 557026 17778 557262 18014
rect 556706 -4422 556942 -4186
rect 557026 -4422 557262 -4186
rect 556706 -4742 556942 -4506
rect 557026 -4742 557262 -4506
rect 560426 709402 560662 709638
rect 560746 709402 560982 709638
rect 560426 709082 560662 709318
rect 560746 709082 560982 709318
rect 560426 669818 560662 670054
rect 560746 669818 560982 670054
rect 560426 669498 560662 669734
rect 560746 669498 560982 669734
rect 560426 633818 560662 634054
rect 560746 633818 560982 634054
rect 560426 633498 560662 633734
rect 560746 633498 560982 633734
rect 560426 597818 560662 598054
rect 560746 597818 560982 598054
rect 560426 597498 560662 597734
rect 560746 597498 560982 597734
rect 560426 561818 560662 562054
rect 560746 561818 560982 562054
rect 560426 561498 560662 561734
rect 560746 561498 560982 561734
rect 560426 525818 560662 526054
rect 560746 525818 560982 526054
rect 560426 525498 560662 525734
rect 560746 525498 560982 525734
rect 560426 489818 560662 490054
rect 560746 489818 560982 490054
rect 560426 489498 560662 489734
rect 560746 489498 560982 489734
rect 560426 453818 560662 454054
rect 560746 453818 560982 454054
rect 560426 453498 560662 453734
rect 560746 453498 560982 453734
rect 560426 417818 560662 418054
rect 560746 417818 560982 418054
rect 560426 417498 560662 417734
rect 560746 417498 560982 417734
rect 560426 381818 560662 382054
rect 560746 381818 560982 382054
rect 560426 381498 560662 381734
rect 560746 381498 560982 381734
rect 560426 345818 560662 346054
rect 560746 345818 560982 346054
rect 560426 345498 560662 345734
rect 560746 345498 560982 345734
rect 560426 309818 560662 310054
rect 560746 309818 560982 310054
rect 560426 309498 560662 309734
rect 560746 309498 560982 309734
rect 560426 273818 560662 274054
rect 560746 273818 560982 274054
rect 560426 273498 560662 273734
rect 560746 273498 560982 273734
rect 560426 237818 560662 238054
rect 560746 237818 560982 238054
rect 560426 237498 560662 237734
rect 560746 237498 560982 237734
rect 560426 201818 560662 202054
rect 560746 201818 560982 202054
rect 560426 201498 560662 201734
rect 560746 201498 560982 201734
rect 560426 165818 560662 166054
rect 560746 165818 560982 166054
rect 560426 165498 560662 165734
rect 560746 165498 560982 165734
rect 560426 129818 560662 130054
rect 560746 129818 560982 130054
rect 560426 129498 560662 129734
rect 560746 129498 560982 129734
rect 560426 93818 560662 94054
rect 560746 93818 560982 94054
rect 560426 93498 560662 93734
rect 560746 93498 560982 93734
rect 560426 57818 560662 58054
rect 560746 57818 560982 58054
rect 560426 57498 560662 57734
rect 560746 57498 560982 57734
rect 560426 21818 560662 22054
rect 560746 21818 560982 22054
rect 560426 21498 560662 21734
rect 560746 21498 560982 21734
rect 560426 -5382 560662 -5146
rect 560746 -5382 560982 -5146
rect 560426 -5702 560662 -5466
rect 560746 -5702 560982 -5466
rect 564146 710362 564382 710598
rect 564466 710362 564702 710598
rect 564146 710042 564382 710278
rect 564466 710042 564702 710278
rect 564146 673538 564382 673774
rect 564466 673538 564702 673774
rect 564146 673218 564382 673454
rect 564466 673218 564702 673454
rect 564146 637538 564382 637774
rect 564466 637538 564702 637774
rect 564146 637218 564382 637454
rect 564466 637218 564702 637454
rect 564146 601538 564382 601774
rect 564466 601538 564702 601774
rect 564146 601218 564382 601454
rect 564466 601218 564702 601454
rect 564146 565538 564382 565774
rect 564466 565538 564702 565774
rect 564146 565218 564382 565454
rect 564466 565218 564702 565454
rect 564146 529538 564382 529774
rect 564466 529538 564702 529774
rect 564146 529218 564382 529454
rect 564466 529218 564702 529454
rect 564146 493538 564382 493774
rect 564466 493538 564702 493774
rect 564146 493218 564382 493454
rect 564466 493218 564702 493454
rect 564146 457538 564382 457774
rect 564466 457538 564702 457774
rect 564146 457218 564382 457454
rect 564466 457218 564702 457454
rect 564146 421538 564382 421774
rect 564466 421538 564702 421774
rect 564146 421218 564382 421454
rect 564466 421218 564702 421454
rect 564146 385538 564382 385774
rect 564466 385538 564702 385774
rect 564146 385218 564382 385454
rect 564466 385218 564702 385454
rect 564146 349538 564382 349774
rect 564466 349538 564702 349774
rect 564146 349218 564382 349454
rect 564466 349218 564702 349454
rect 564146 313538 564382 313774
rect 564466 313538 564702 313774
rect 564146 313218 564382 313454
rect 564466 313218 564702 313454
rect 564146 277538 564382 277774
rect 564466 277538 564702 277774
rect 564146 277218 564382 277454
rect 564466 277218 564702 277454
rect 564146 241538 564382 241774
rect 564466 241538 564702 241774
rect 564146 241218 564382 241454
rect 564466 241218 564702 241454
rect 564146 205538 564382 205774
rect 564466 205538 564702 205774
rect 564146 205218 564382 205454
rect 564466 205218 564702 205454
rect 564146 169538 564382 169774
rect 564466 169538 564702 169774
rect 564146 169218 564382 169454
rect 564466 169218 564702 169454
rect 564146 133538 564382 133774
rect 564466 133538 564702 133774
rect 564146 133218 564382 133454
rect 564466 133218 564702 133454
rect 564146 97538 564382 97774
rect 564466 97538 564702 97774
rect 564146 97218 564382 97454
rect 564466 97218 564702 97454
rect 564146 61538 564382 61774
rect 564466 61538 564702 61774
rect 564146 61218 564382 61454
rect 564466 61218 564702 61454
rect 564146 25538 564382 25774
rect 564466 25538 564702 25774
rect 564146 25218 564382 25454
rect 564466 25218 564702 25454
rect 564146 -6342 564382 -6106
rect 564466 -6342 564702 -6106
rect 564146 -6662 564382 -6426
rect 564466 -6662 564702 -6426
rect 567866 711322 568102 711558
rect 568186 711322 568422 711558
rect 567866 711002 568102 711238
rect 568186 711002 568422 711238
rect 567866 677258 568102 677494
rect 568186 677258 568422 677494
rect 567866 676938 568102 677174
rect 568186 676938 568422 677174
rect 567866 641258 568102 641494
rect 568186 641258 568422 641494
rect 567866 640938 568102 641174
rect 568186 640938 568422 641174
rect 567866 605258 568102 605494
rect 568186 605258 568422 605494
rect 567866 604938 568102 605174
rect 568186 604938 568422 605174
rect 567866 569258 568102 569494
rect 568186 569258 568422 569494
rect 567866 568938 568102 569174
rect 568186 568938 568422 569174
rect 567866 533258 568102 533494
rect 568186 533258 568422 533494
rect 567866 532938 568102 533174
rect 568186 532938 568422 533174
rect 567866 497258 568102 497494
rect 568186 497258 568422 497494
rect 567866 496938 568102 497174
rect 568186 496938 568422 497174
rect 567866 461258 568102 461494
rect 568186 461258 568422 461494
rect 567866 460938 568102 461174
rect 568186 460938 568422 461174
rect 567866 425258 568102 425494
rect 568186 425258 568422 425494
rect 567866 424938 568102 425174
rect 568186 424938 568422 425174
rect 567866 389258 568102 389494
rect 568186 389258 568422 389494
rect 567866 388938 568102 389174
rect 568186 388938 568422 389174
rect 567866 353258 568102 353494
rect 568186 353258 568422 353494
rect 567866 352938 568102 353174
rect 568186 352938 568422 353174
rect 567866 317258 568102 317494
rect 568186 317258 568422 317494
rect 567866 316938 568102 317174
rect 568186 316938 568422 317174
rect 567866 281258 568102 281494
rect 568186 281258 568422 281494
rect 567866 280938 568102 281174
rect 568186 280938 568422 281174
rect 567866 245258 568102 245494
rect 568186 245258 568422 245494
rect 567866 244938 568102 245174
rect 568186 244938 568422 245174
rect 567866 209258 568102 209494
rect 568186 209258 568422 209494
rect 567866 208938 568102 209174
rect 568186 208938 568422 209174
rect 567866 173258 568102 173494
rect 568186 173258 568422 173494
rect 567866 172938 568102 173174
rect 568186 172938 568422 173174
rect 567866 137258 568102 137494
rect 568186 137258 568422 137494
rect 567866 136938 568102 137174
rect 568186 136938 568422 137174
rect 567866 101258 568102 101494
rect 568186 101258 568422 101494
rect 567866 100938 568102 101174
rect 568186 100938 568422 101174
rect 567866 65258 568102 65494
rect 568186 65258 568422 65494
rect 567866 64938 568102 65174
rect 568186 64938 568422 65174
rect 567866 29258 568102 29494
rect 568186 29258 568422 29494
rect 567866 28938 568102 29174
rect 568186 28938 568422 29174
rect 567866 -7302 568102 -7066
rect 568186 -7302 568422 -7066
rect 567866 -7622 568102 -7386
rect 568186 -7622 568422 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 690938 586538 691174
rect 586622 690938 586858 691174
rect 586302 690618 586538 690854
rect 586622 690618 586858 690854
rect 586302 654938 586538 655174
rect 586622 654938 586858 655174
rect 586302 654618 586538 654854
rect 586622 654618 586858 654854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 582938 586538 583174
rect 586622 582938 586858 583174
rect 586302 582618 586538 582854
rect 586622 582618 586858 582854
rect 586302 546938 586538 547174
rect 586622 546938 586858 547174
rect 586302 546618 586538 546854
rect 586622 546618 586858 546854
rect 586302 510938 586538 511174
rect 586622 510938 586858 511174
rect 586302 510618 586538 510854
rect 586622 510618 586858 510854
rect 586302 474938 586538 475174
rect 586622 474938 586858 475174
rect 586302 474618 586538 474854
rect 586622 474618 586858 474854
rect 586302 438938 586538 439174
rect 586622 438938 586858 439174
rect 586302 438618 586538 438854
rect 586622 438618 586858 438854
rect 586302 402938 586538 403174
rect 586622 402938 586858 403174
rect 586302 402618 586538 402854
rect 586622 402618 586858 402854
rect 586302 366938 586538 367174
rect 586622 366938 586858 367174
rect 586302 366618 586538 366854
rect 586622 366618 586858 366854
rect 586302 330938 586538 331174
rect 586622 330938 586858 331174
rect 586302 330618 586538 330854
rect 586622 330618 586858 330854
rect 586302 294938 586538 295174
rect 586622 294938 586858 295174
rect 586302 294618 586538 294854
rect 586622 294618 586858 294854
rect 586302 258938 586538 259174
rect 586622 258938 586858 259174
rect 586302 258618 586538 258854
rect 586622 258618 586858 258854
rect 586302 222938 586538 223174
rect 586622 222938 586858 223174
rect 586302 222618 586538 222854
rect 586622 222618 586858 222854
rect 586302 186938 586538 187174
rect 586622 186938 586858 187174
rect 586302 186618 586538 186854
rect 586622 186618 586858 186854
rect 586302 150938 586538 151174
rect 586622 150938 586858 151174
rect 586302 150618 586538 150854
rect 586622 150618 586858 150854
rect 586302 114938 586538 115174
rect 586622 114938 586858 115174
rect 586302 114618 586538 114854
rect 586622 114618 586858 114854
rect 586302 78938 586538 79174
rect 586622 78938 586858 79174
rect 586302 78618 586538 78854
rect 586622 78618 586858 78854
rect 586302 42938 586538 43174
rect 586622 42938 586858 43174
rect 586302 42618 586538 42854
rect 586622 42618 586858 42854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 694658 587498 694894
rect 587582 694658 587818 694894
rect 587262 694338 587498 694574
rect 587582 694338 587818 694574
rect 587262 658658 587498 658894
rect 587582 658658 587818 658894
rect 587262 658338 587498 658574
rect 587582 658338 587818 658574
rect 587262 622658 587498 622894
rect 587582 622658 587818 622894
rect 587262 622338 587498 622574
rect 587582 622338 587818 622574
rect 587262 586658 587498 586894
rect 587582 586658 587818 586894
rect 587262 586338 587498 586574
rect 587582 586338 587818 586574
rect 587262 550658 587498 550894
rect 587582 550658 587818 550894
rect 587262 550338 587498 550574
rect 587582 550338 587818 550574
rect 587262 514658 587498 514894
rect 587582 514658 587818 514894
rect 587262 514338 587498 514574
rect 587582 514338 587818 514574
rect 587262 478658 587498 478894
rect 587582 478658 587818 478894
rect 587262 478338 587498 478574
rect 587582 478338 587818 478574
rect 587262 442658 587498 442894
rect 587582 442658 587818 442894
rect 587262 442338 587498 442574
rect 587582 442338 587818 442574
rect 587262 406658 587498 406894
rect 587582 406658 587818 406894
rect 587262 406338 587498 406574
rect 587582 406338 587818 406574
rect 587262 370658 587498 370894
rect 587582 370658 587818 370894
rect 587262 370338 587498 370574
rect 587582 370338 587818 370574
rect 587262 334658 587498 334894
rect 587582 334658 587818 334894
rect 587262 334338 587498 334574
rect 587582 334338 587818 334574
rect 587262 298658 587498 298894
rect 587582 298658 587818 298894
rect 587262 298338 587498 298574
rect 587582 298338 587818 298574
rect 587262 262658 587498 262894
rect 587582 262658 587818 262894
rect 587262 262338 587498 262574
rect 587582 262338 587818 262574
rect 587262 226658 587498 226894
rect 587582 226658 587818 226894
rect 587262 226338 587498 226574
rect 587582 226338 587818 226574
rect 587262 190658 587498 190894
rect 587582 190658 587818 190894
rect 587262 190338 587498 190574
rect 587582 190338 587818 190574
rect 587262 154658 587498 154894
rect 587582 154658 587818 154894
rect 587262 154338 587498 154574
rect 587582 154338 587818 154574
rect 587262 118658 587498 118894
rect 587582 118658 587818 118894
rect 587262 118338 587498 118574
rect 587582 118338 587818 118574
rect 587262 82658 587498 82894
rect 587582 82658 587818 82894
rect 587262 82338 587498 82574
rect 587582 82338 587818 82574
rect 587262 46658 587498 46894
rect 587582 46658 587818 46894
rect 587262 46338 587498 46574
rect 587582 46338 587818 46574
rect 587262 10658 587498 10894
rect 587582 10658 587818 10894
rect 587262 10338 587498 10574
rect 587582 10338 587818 10574
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 698378 588458 698614
rect 588542 698378 588778 698614
rect 588222 698058 588458 698294
rect 588542 698058 588778 698294
rect 588222 662378 588458 662614
rect 588542 662378 588778 662614
rect 588222 662058 588458 662294
rect 588542 662058 588778 662294
rect 588222 626378 588458 626614
rect 588542 626378 588778 626614
rect 588222 626058 588458 626294
rect 588542 626058 588778 626294
rect 588222 590378 588458 590614
rect 588542 590378 588778 590614
rect 588222 590058 588458 590294
rect 588542 590058 588778 590294
rect 588222 554378 588458 554614
rect 588542 554378 588778 554614
rect 588222 554058 588458 554294
rect 588542 554058 588778 554294
rect 588222 518378 588458 518614
rect 588542 518378 588778 518614
rect 588222 518058 588458 518294
rect 588542 518058 588778 518294
rect 588222 482378 588458 482614
rect 588542 482378 588778 482614
rect 588222 482058 588458 482294
rect 588542 482058 588778 482294
rect 588222 446378 588458 446614
rect 588542 446378 588778 446614
rect 588222 446058 588458 446294
rect 588542 446058 588778 446294
rect 588222 410378 588458 410614
rect 588542 410378 588778 410614
rect 588222 410058 588458 410294
rect 588542 410058 588778 410294
rect 588222 374378 588458 374614
rect 588542 374378 588778 374614
rect 588222 374058 588458 374294
rect 588542 374058 588778 374294
rect 588222 338378 588458 338614
rect 588542 338378 588778 338614
rect 588222 338058 588458 338294
rect 588542 338058 588778 338294
rect 588222 302378 588458 302614
rect 588542 302378 588778 302614
rect 588222 302058 588458 302294
rect 588542 302058 588778 302294
rect 588222 266378 588458 266614
rect 588542 266378 588778 266614
rect 588222 266058 588458 266294
rect 588542 266058 588778 266294
rect 588222 230378 588458 230614
rect 588542 230378 588778 230614
rect 588222 230058 588458 230294
rect 588542 230058 588778 230294
rect 588222 194378 588458 194614
rect 588542 194378 588778 194614
rect 588222 194058 588458 194294
rect 588542 194058 588778 194294
rect 588222 158378 588458 158614
rect 588542 158378 588778 158614
rect 588222 158058 588458 158294
rect 588542 158058 588778 158294
rect 588222 122378 588458 122614
rect 588542 122378 588778 122614
rect 588222 122058 588458 122294
rect 588542 122058 588778 122294
rect 588222 86378 588458 86614
rect 588542 86378 588778 86614
rect 588222 86058 588458 86294
rect 588542 86058 588778 86294
rect 588222 50378 588458 50614
rect 588542 50378 588778 50614
rect 588222 50058 588458 50294
rect 588542 50058 588778 50294
rect 588222 14378 588458 14614
rect 588542 14378 588778 14614
rect 588222 14058 588458 14294
rect 588542 14058 588778 14294
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 666098 589418 666334
rect 589502 666098 589738 666334
rect 589182 665778 589418 666014
rect 589502 665778 589738 666014
rect 589182 630098 589418 630334
rect 589502 630098 589738 630334
rect 589182 629778 589418 630014
rect 589502 629778 589738 630014
rect 589182 594098 589418 594334
rect 589502 594098 589738 594334
rect 589182 593778 589418 594014
rect 589502 593778 589738 594014
rect 589182 558098 589418 558334
rect 589502 558098 589738 558334
rect 589182 557778 589418 558014
rect 589502 557778 589738 558014
rect 589182 522098 589418 522334
rect 589502 522098 589738 522334
rect 589182 521778 589418 522014
rect 589502 521778 589738 522014
rect 589182 486098 589418 486334
rect 589502 486098 589738 486334
rect 589182 485778 589418 486014
rect 589502 485778 589738 486014
rect 589182 450098 589418 450334
rect 589502 450098 589738 450334
rect 589182 449778 589418 450014
rect 589502 449778 589738 450014
rect 589182 414098 589418 414334
rect 589502 414098 589738 414334
rect 589182 413778 589418 414014
rect 589502 413778 589738 414014
rect 589182 378098 589418 378334
rect 589502 378098 589738 378334
rect 589182 377778 589418 378014
rect 589502 377778 589738 378014
rect 589182 342098 589418 342334
rect 589502 342098 589738 342334
rect 589182 341778 589418 342014
rect 589502 341778 589738 342014
rect 589182 306098 589418 306334
rect 589502 306098 589738 306334
rect 589182 305778 589418 306014
rect 589502 305778 589738 306014
rect 589182 270098 589418 270334
rect 589502 270098 589738 270334
rect 589182 269778 589418 270014
rect 589502 269778 589738 270014
rect 589182 234098 589418 234334
rect 589502 234098 589738 234334
rect 589182 233778 589418 234014
rect 589502 233778 589738 234014
rect 589182 198098 589418 198334
rect 589502 198098 589738 198334
rect 589182 197778 589418 198014
rect 589502 197778 589738 198014
rect 589182 162098 589418 162334
rect 589502 162098 589738 162334
rect 589182 161778 589418 162014
rect 589502 161778 589738 162014
rect 589182 126098 589418 126334
rect 589502 126098 589738 126334
rect 589182 125778 589418 126014
rect 589502 125778 589738 126014
rect 589182 90098 589418 90334
rect 589502 90098 589738 90334
rect 589182 89778 589418 90014
rect 589502 89778 589738 90014
rect 589182 54098 589418 54334
rect 589502 54098 589738 54334
rect 589182 53778 589418 54014
rect 589502 53778 589738 54014
rect 589182 18098 589418 18334
rect 589502 18098 589738 18334
rect 589182 17778 589418 18014
rect 589502 17778 589738 18014
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 669818 590378 670054
rect 590462 669818 590698 670054
rect 590142 669498 590378 669734
rect 590462 669498 590698 669734
rect 590142 633818 590378 634054
rect 590462 633818 590698 634054
rect 590142 633498 590378 633734
rect 590462 633498 590698 633734
rect 590142 597818 590378 598054
rect 590462 597818 590698 598054
rect 590142 597498 590378 597734
rect 590462 597498 590698 597734
rect 590142 561818 590378 562054
rect 590462 561818 590698 562054
rect 590142 561498 590378 561734
rect 590462 561498 590698 561734
rect 590142 525818 590378 526054
rect 590462 525818 590698 526054
rect 590142 525498 590378 525734
rect 590462 525498 590698 525734
rect 590142 489818 590378 490054
rect 590462 489818 590698 490054
rect 590142 489498 590378 489734
rect 590462 489498 590698 489734
rect 590142 453818 590378 454054
rect 590462 453818 590698 454054
rect 590142 453498 590378 453734
rect 590462 453498 590698 453734
rect 590142 417818 590378 418054
rect 590462 417818 590698 418054
rect 590142 417498 590378 417734
rect 590462 417498 590698 417734
rect 590142 381818 590378 382054
rect 590462 381818 590698 382054
rect 590142 381498 590378 381734
rect 590462 381498 590698 381734
rect 590142 345818 590378 346054
rect 590462 345818 590698 346054
rect 590142 345498 590378 345734
rect 590462 345498 590698 345734
rect 590142 309818 590378 310054
rect 590462 309818 590698 310054
rect 590142 309498 590378 309734
rect 590462 309498 590698 309734
rect 590142 273818 590378 274054
rect 590462 273818 590698 274054
rect 590142 273498 590378 273734
rect 590462 273498 590698 273734
rect 590142 237818 590378 238054
rect 590462 237818 590698 238054
rect 590142 237498 590378 237734
rect 590462 237498 590698 237734
rect 590142 201818 590378 202054
rect 590462 201818 590698 202054
rect 590142 201498 590378 201734
rect 590462 201498 590698 201734
rect 590142 165818 590378 166054
rect 590462 165818 590698 166054
rect 590142 165498 590378 165734
rect 590462 165498 590698 165734
rect 590142 129818 590378 130054
rect 590462 129818 590698 130054
rect 590142 129498 590378 129734
rect 590462 129498 590698 129734
rect 590142 93818 590378 94054
rect 590462 93818 590698 94054
rect 590142 93498 590378 93734
rect 590462 93498 590698 93734
rect 590142 57818 590378 58054
rect 590462 57818 590698 58054
rect 590142 57498 590378 57734
rect 590462 57498 590698 57734
rect 590142 21818 590378 22054
rect 590462 21818 590698 22054
rect 590142 21498 590378 21734
rect 590462 21498 590698 21734
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 673538 591338 673774
rect 591422 673538 591658 673774
rect 591102 673218 591338 673454
rect 591422 673218 591658 673454
rect 591102 637538 591338 637774
rect 591422 637538 591658 637774
rect 591102 637218 591338 637454
rect 591422 637218 591658 637454
rect 591102 601538 591338 601774
rect 591422 601538 591658 601774
rect 591102 601218 591338 601454
rect 591422 601218 591658 601454
rect 591102 565538 591338 565774
rect 591422 565538 591658 565774
rect 591102 565218 591338 565454
rect 591422 565218 591658 565454
rect 591102 529538 591338 529774
rect 591422 529538 591658 529774
rect 591102 529218 591338 529454
rect 591422 529218 591658 529454
rect 591102 493538 591338 493774
rect 591422 493538 591658 493774
rect 591102 493218 591338 493454
rect 591422 493218 591658 493454
rect 591102 457538 591338 457774
rect 591422 457538 591658 457774
rect 591102 457218 591338 457454
rect 591422 457218 591658 457454
rect 591102 421538 591338 421774
rect 591422 421538 591658 421774
rect 591102 421218 591338 421454
rect 591422 421218 591658 421454
rect 591102 385538 591338 385774
rect 591422 385538 591658 385774
rect 591102 385218 591338 385454
rect 591422 385218 591658 385454
rect 591102 349538 591338 349774
rect 591422 349538 591658 349774
rect 591102 349218 591338 349454
rect 591422 349218 591658 349454
rect 591102 313538 591338 313774
rect 591422 313538 591658 313774
rect 591102 313218 591338 313454
rect 591422 313218 591658 313454
rect 591102 277538 591338 277774
rect 591422 277538 591658 277774
rect 591102 277218 591338 277454
rect 591422 277218 591658 277454
rect 591102 241538 591338 241774
rect 591422 241538 591658 241774
rect 591102 241218 591338 241454
rect 591422 241218 591658 241454
rect 591102 205538 591338 205774
rect 591422 205538 591658 205774
rect 591102 205218 591338 205454
rect 591422 205218 591658 205454
rect 591102 169538 591338 169774
rect 591422 169538 591658 169774
rect 591102 169218 591338 169454
rect 591422 169218 591658 169454
rect 591102 133538 591338 133774
rect 591422 133538 591658 133774
rect 591102 133218 591338 133454
rect 591422 133218 591658 133454
rect 591102 97538 591338 97774
rect 591422 97538 591658 97774
rect 591102 97218 591338 97454
rect 591422 97218 591658 97454
rect 591102 61538 591338 61774
rect 591422 61538 591658 61774
rect 591102 61218 591338 61454
rect 591422 61218 591658 61454
rect 591102 25538 591338 25774
rect 591422 25538 591658 25774
rect 591102 25218 591338 25454
rect 591422 25218 591658 25454
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 677258 592298 677494
rect 592382 677258 592618 677494
rect 592062 676938 592298 677174
rect 592382 676938 592618 677174
rect 592062 641258 592298 641494
rect 592382 641258 592618 641494
rect 592062 640938 592298 641174
rect 592382 640938 592618 641174
rect 592062 605258 592298 605494
rect 592382 605258 592618 605494
rect 592062 604938 592298 605174
rect 592382 604938 592618 605174
rect 592062 569258 592298 569494
rect 592382 569258 592618 569494
rect 592062 568938 592298 569174
rect 592382 568938 592618 569174
rect 592062 533258 592298 533494
rect 592382 533258 592618 533494
rect 592062 532938 592298 533174
rect 592382 532938 592618 533174
rect 592062 497258 592298 497494
rect 592382 497258 592618 497494
rect 592062 496938 592298 497174
rect 592382 496938 592618 497174
rect 592062 461258 592298 461494
rect 592382 461258 592618 461494
rect 592062 460938 592298 461174
rect 592382 460938 592618 461174
rect 592062 425258 592298 425494
rect 592382 425258 592618 425494
rect 592062 424938 592298 425174
rect 592382 424938 592618 425174
rect 592062 389258 592298 389494
rect 592382 389258 592618 389494
rect 592062 388938 592298 389174
rect 592382 388938 592618 389174
rect 592062 353258 592298 353494
rect 592382 353258 592618 353494
rect 592062 352938 592298 353174
rect 592382 352938 592618 353174
rect 592062 317258 592298 317494
rect 592382 317258 592618 317494
rect 592062 316938 592298 317174
rect 592382 316938 592618 317174
rect 592062 281258 592298 281494
rect 592382 281258 592618 281494
rect 592062 280938 592298 281174
rect 592382 280938 592618 281174
rect 592062 245258 592298 245494
rect 592382 245258 592618 245494
rect 592062 244938 592298 245174
rect 592382 244938 592618 245174
rect 592062 209258 592298 209494
rect 592382 209258 592618 209494
rect 592062 208938 592298 209174
rect 592382 208938 592618 209174
rect 592062 173258 592298 173494
rect 592382 173258 592618 173494
rect 592062 172938 592298 173174
rect 592382 172938 592618 173174
rect 592062 137258 592298 137494
rect 592382 137258 592618 137494
rect 592062 136938 592298 137174
rect 592382 136938 592618 137174
rect 592062 101258 592298 101494
rect 592382 101258 592618 101494
rect 592062 100938 592298 101174
rect 592382 100938 592618 101174
rect 592062 65258 592298 65494
rect 592382 65258 592618 65494
rect 592062 64938 592298 65174
rect 592382 64938 592618 65174
rect 592062 29258 592298 29494
rect 592382 29258 592618 29494
rect 592062 28938 592298 29174
rect 592382 28938 592618 29174
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 315866 711558
rect 316102 711322 316186 711558
rect 316422 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 315866 711238
rect 316102 711002 316186 711238
rect 316422 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 24146 710598
rect 24382 710362 24466 710598
rect 24702 710362 60146 710598
rect 60382 710362 60466 710598
rect 60702 710362 96146 710598
rect 96382 710362 96466 710598
rect 96702 710362 132146 710598
rect 132382 710362 132466 710598
rect 132702 710362 168146 710598
rect 168382 710362 168466 710598
rect 168702 710362 204146 710598
rect 204382 710362 204466 710598
rect 204702 710362 240146 710598
rect 240382 710362 240466 710598
rect 240702 710362 276146 710598
rect 276382 710362 276466 710598
rect 276702 710362 312146 710598
rect 312382 710362 312466 710598
rect 312702 710362 348146 710598
rect 348382 710362 348466 710598
rect 348702 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 24146 710278
rect 24382 710042 24466 710278
rect 24702 710042 60146 710278
rect 60382 710042 60466 710278
rect 60702 710042 96146 710278
rect 96382 710042 96466 710278
rect 96702 710042 132146 710278
rect 132382 710042 132466 710278
rect 132702 710042 168146 710278
rect 168382 710042 168466 710278
rect 168702 710042 204146 710278
rect 204382 710042 204466 710278
rect 204702 710042 240146 710278
rect 240382 710042 240466 710278
rect 240702 710042 276146 710278
rect 276382 710042 276466 710278
rect 276702 710042 312146 710278
rect 312382 710042 312466 710278
rect 312702 710042 348146 710278
rect 348382 710042 348466 710278
rect 348702 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 56426 709638
rect 56662 709402 56746 709638
rect 56982 709402 92426 709638
rect 92662 709402 92746 709638
rect 92982 709402 128426 709638
rect 128662 709402 128746 709638
rect 128982 709402 164426 709638
rect 164662 709402 164746 709638
rect 164982 709402 200426 709638
rect 200662 709402 200746 709638
rect 200982 709402 236426 709638
rect 236662 709402 236746 709638
rect 236982 709402 272426 709638
rect 272662 709402 272746 709638
rect 272982 709402 308426 709638
rect 308662 709402 308746 709638
rect 308982 709402 344426 709638
rect 344662 709402 344746 709638
rect 344982 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 56426 709318
rect 56662 709082 56746 709318
rect 56982 709082 92426 709318
rect 92662 709082 92746 709318
rect 92982 709082 128426 709318
rect 128662 709082 128746 709318
rect 128982 709082 164426 709318
rect 164662 709082 164746 709318
rect 164982 709082 200426 709318
rect 200662 709082 200746 709318
rect 200982 709082 236426 709318
rect 236662 709082 236746 709318
rect 236982 709082 272426 709318
rect 272662 709082 272746 709318
rect 272982 709082 308426 709318
rect 308662 709082 308746 709318
rect 308982 709082 344426 709318
rect 344662 709082 344746 709318
rect 344982 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 52706 708678
rect 52942 708442 53026 708678
rect 53262 708442 88706 708678
rect 88942 708442 89026 708678
rect 89262 708442 124706 708678
rect 124942 708442 125026 708678
rect 125262 708442 160706 708678
rect 160942 708442 161026 708678
rect 161262 708442 196706 708678
rect 196942 708442 197026 708678
rect 197262 708442 232706 708678
rect 232942 708442 233026 708678
rect 233262 708442 268706 708678
rect 268942 708442 269026 708678
rect 269262 708442 304706 708678
rect 304942 708442 305026 708678
rect 305262 708442 340706 708678
rect 340942 708442 341026 708678
rect 341262 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 484706 708678
rect 484942 708442 485026 708678
rect 485262 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 52706 708358
rect 52942 708122 53026 708358
rect 53262 708122 88706 708358
rect 88942 708122 89026 708358
rect 89262 708122 124706 708358
rect 124942 708122 125026 708358
rect 125262 708122 160706 708358
rect 160942 708122 161026 708358
rect 161262 708122 196706 708358
rect 196942 708122 197026 708358
rect 197262 708122 232706 708358
rect 232942 708122 233026 708358
rect 233262 708122 268706 708358
rect 268942 708122 269026 708358
rect 269262 708122 304706 708358
rect 304942 708122 305026 708358
rect 305262 708122 340706 708358
rect 340942 708122 341026 708358
rect 341262 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 484706 708358
rect 484942 708122 485026 708358
rect 485262 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 592650 698294
rect -8726 698026 592650 698058
rect -8726 694894 592650 694926
rect -8726 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 592650 694894
rect -8726 694574 592650 694658
rect -8726 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 592650 694574
rect -8726 694306 592650 694338
rect -8726 691174 592650 691206
rect -8726 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 592650 691174
rect -8726 690854 592650 690938
rect -8726 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 592650 690854
rect -8726 690586 592650 690618
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 677494 592650 677526
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 315866 677494
rect 316102 677258 316186 677494
rect 316422 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect -8726 677174 592650 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 315866 677174
rect 316102 676938 316186 677174
rect 316422 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect -8726 676906 592650 676938
rect -8726 673774 592650 673806
rect -8726 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 24146 673774
rect 24382 673538 24466 673774
rect 24702 673538 60146 673774
rect 60382 673538 60466 673774
rect 60702 673538 96146 673774
rect 96382 673538 96466 673774
rect 96702 673538 132146 673774
rect 132382 673538 132466 673774
rect 132702 673538 168146 673774
rect 168382 673538 168466 673774
rect 168702 673538 204146 673774
rect 204382 673538 204466 673774
rect 204702 673538 240146 673774
rect 240382 673538 240466 673774
rect 240702 673538 276146 673774
rect 276382 673538 276466 673774
rect 276702 673538 312146 673774
rect 312382 673538 312466 673774
rect 312702 673538 348146 673774
rect 348382 673538 348466 673774
rect 348702 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 592650 673774
rect -8726 673454 592650 673538
rect -8726 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 24146 673454
rect 24382 673218 24466 673454
rect 24702 673218 60146 673454
rect 60382 673218 60466 673454
rect 60702 673218 96146 673454
rect 96382 673218 96466 673454
rect 96702 673218 132146 673454
rect 132382 673218 132466 673454
rect 132702 673218 168146 673454
rect 168382 673218 168466 673454
rect 168702 673218 204146 673454
rect 204382 673218 204466 673454
rect 204702 673218 240146 673454
rect 240382 673218 240466 673454
rect 240702 673218 276146 673454
rect 276382 673218 276466 673454
rect 276702 673218 312146 673454
rect 312382 673218 312466 673454
rect 312702 673218 348146 673454
rect 348382 673218 348466 673454
rect 348702 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 592650 673454
rect -8726 673186 592650 673218
rect -8726 670054 592650 670086
rect -8726 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 56426 670054
rect 56662 669818 56746 670054
rect 56982 669818 92426 670054
rect 92662 669818 92746 670054
rect 92982 669818 128426 670054
rect 128662 669818 128746 670054
rect 128982 669818 164426 670054
rect 164662 669818 164746 670054
rect 164982 669818 200426 670054
rect 200662 669818 200746 670054
rect 200982 669818 236426 670054
rect 236662 669818 236746 670054
rect 236982 669818 272426 670054
rect 272662 669818 272746 670054
rect 272982 669818 308426 670054
rect 308662 669818 308746 670054
rect 308982 669818 344426 670054
rect 344662 669818 344746 670054
rect 344982 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 592650 670054
rect -8726 669734 592650 669818
rect -8726 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 56426 669734
rect 56662 669498 56746 669734
rect 56982 669498 92426 669734
rect 92662 669498 92746 669734
rect 92982 669498 128426 669734
rect 128662 669498 128746 669734
rect 128982 669498 164426 669734
rect 164662 669498 164746 669734
rect 164982 669498 200426 669734
rect 200662 669498 200746 669734
rect 200982 669498 236426 669734
rect 236662 669498 236746 669734
rect 236982 669498 272426 669734
rect 272662 669498 272746 669734
rect 272982 669498 308426 669734
rect 308662 669498 308746 669734
rect 308982 669498 344426 669734
rect 344662 669498 344746 669734
rect 344982 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 592650 669734
rect -8726 669466 592650 669498
rect -8726 666334 592650 666366
rect -8726 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 52706 666334
rect 52942 666098 53026 666334
rect 53262 666098 88706 666334
rect 88942 666098 89026 666334
rect 89262 666098 124706 666334
rect 124942 666098 125026 666334
rect 125262 666098 160706 666334
rect 160942 666098 161026 666334
rect 161262 666098 196706 666334
rect 196942 666098 197026 666334
rect 197262 666098 232706 666334
rect 232942 666098 233026 666334
rect 233262 666098 268706 666334
rect 268942 666098 269026 666334
rect 269262 666098 304706 666334
rect 304942 666098 305026 666334
rect 305262 666098 340706 666334
rect 340942 666098 341026 666334
rect 341262 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 484706 666334
rect 484942 666098 485026 666334
rect 485262 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 592650 666334
rect -8726 666014 592650 666098
rect -8726 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 52706 666014
rect 52942 665778 53026 666014
rect 53262 665778 88706 666014
rect 88942 665778 89026 666014
rect 89262 665778 124706 666014
rect 124942 665778 125026 666014
rect 125262 665778 160706 666014
rect 160942 665778 161026 666014
rect 161262 665778 196706 666014
rect 196942 665778 197026 666014
rect 197262 665778 232706 666014
rect 232942 665778 233026 666014
rect 233262 665778 268706 666014
rect 268942 665778 269026 666014
rect 269262 665778 304706 666014
rect 304942 665778 305026 666014
rect 305262 665778 340706 666014
rect 340942 665778 341026 666014
rect 341262 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 484706 666014
rect 484942 665778 485026 666014
rect 485262 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 592650 666014
rect -8726 665746 592650 665778
rect -8726 662614 592650 662646
rect -8726 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 592650 662294
rect -8726 662026 592650 662058
rect -8726 658894 592650 658926
rect -8726 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 592650 658894
rect -8726 658574 592650 658658
rect -8726 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 592650 658574
rect -8726 658306 592650 658338
rect -8726 655174 592650 655206
rect -8726 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 592650 655174
rect -8726 654854 592650 654938
rect -8726 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 592650 654854
rect -8726 654586 592650 654618
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 641494 592650 641526
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 63866 641494
rect 64102 641258 64186 641494
rect 64422 641258 99866 641494
rect 100102 641258 100186 641494
rect 100422 641258 135866 641494
rect 136102 641258 136186 641494
rect 136422 641258 171866 641494
rect 172102 641258 172186 641494
rect 172422 641258 207866 641494
rect 208102 641258 208186 641494
rect 208422 641258 243866 641494
rect 244102 641258 244186 641494
rect 244422 641258 279866 641494
rect 280102 641258 280186 641494
rect 280422 641258 315866 641494
rect 316102 641258 316186 641494
rect 316422 641258 351866 641494
rect 352102 641258 352186 641494
rect 352422 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 459866 641494
rect 460102 641258 460186 641494
rect 460422 641258 495866 641494
rect 496102 641258 496186 641494
rect 496422 641258 531866 641494
rect 532102 641258 532186 641494
rect 532422 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect -8726 641174 592650 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 63866 641174
rect 64102 640938 64186 641174
rect 64422 640938 99866 641174
rect 100102 640938 100186 641174
rect 100422 640938 135866 641174
rect 136102 640938 136186 641174
rect 136422 640938 171866 641174
rect 172102 640938 172186 641174
rect 172422 640938 207866 641174
rect 208102 640938 208186 641174
rect 208422 640938 243866 641174
rect 244102 640938 244186 641174
rect 244422 640938 279866 641174
rect 280102 640938 280186 641174
rect 280422 640938 315866 641174
rect 316102 640938 316186 641174
rect 316422 640938 351866 641174
rect 352102 640938 352186 641174
rect 352422 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 459866 641174
rect 460102 640938 460186 641174
rect 460422 640938 495866 641174
rect 496102 640938 496186 641174
rect 496422 640938 531866 641174
rect 532102 640938 532186 641174
rect 532422 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 24146 637774
rect 24382 637538 24466 637774
rect 24702 637538 60146 637774
rect 60382 637538 60466 637774
rect 60702 637538 96146 637774
rect 96382 637538 96466 637774
rect 96702 637538 132146 637774
rect 132382 637538 132466 637774
rect 132702 637538 168146 637774
rect 168382 637538 168466 637774
rect 168702 637538 204146 637774
rect 204382 637538 204466 637774
rect 204702 637538 240146 637774
rect 240382 637538 240466 637774
rect 240702 637538 276146 637774
rect 276382 637538 276466 637774
rect 276702 637538 312146 637774
rect 312382 637538 312466 637774
rect 312702 637538 348146 637774
rect 348382 637538 348466 637774
rect 348702 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 492146 637774
rect 492382 637538 492466 637774
rect 492702 637538 528146 637774
rect 528382 637538 528466 637774
rect 528702 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 592650 637774
rect -8726 637454 592650 637538
rect -8726 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 24146 637454
rect 24382 637218 24466 637454
rect 24702 637218 60146 637454
rect 60382 637218 60466 637454
rect 60702 637218 96146 637454
rect 96382 637218 96466 637454
rect 96702 637218 132146 637454
rect 132382 637218 132466 637454
rect 132702 637218 168146 637454
rect 168382 637218 168466 637454
rect 168702 637218 204146 637454
rect 204382 637218 204466 637454
rect 204702 637218 240146 637454
rect 240382 637218 240466 637454
rect 240702 637218 276146 637454
rect 276382 637218 276466 637454
rect 276702 637218 312146 637454
rect 312382 637218 312466 637454
rect 312702 637218 348146 637454
rect 348382 637218 348466 637454
rect 348702 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 492146 637454
rect 492382 637218 492466 637454
rect 492702 637218 528146 637454
rect 528382 637218 528466 637454
rect 528702 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 592650 637454
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 56426 634054
rect 56662 633818 56746 634054
rect 56982 633818 92426 634054
rect 92662 633818 92746 634054
rect 92982 633818 128426 634054
rect 128662 633818 128746 634054
rect 128982 633818 164426 634054
rect 164662 633818 164746 634054
rect 164982 633818 200426 634054
rect 200662 633818 200746 634054
rect 200982 633818 236426 634054
rect 236662 633818 236746 634054
rect 236982 633818 272426 634054
rect 272662 633818 272746 634054
rect 272982 633818 308426 634054
rect 308662 633818 308746 634054
rect 308982 633818 344426 634054
rect 344662 633818 344746 634054
rect 344982 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 488426 634054
rect 488662 633818 488746 634054
rect 488982 633818 524426 634054
rect 524662 633818 524746 634054
rect 524982 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 592650 634054
rect -8726 633734 592650 633818
rect -8726 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 56426 633734
rect 56662 633498 56746 633734
rect 56982 633498 92426 633734
rect 92662 633498 92746 633734
rect 92982 633498 128426 633734
rect 128662 633498 128746 633734
rect 128982 633498 164426 633734
rect 164662 633498 164746 633734
rect 164982 633498 200426 633734
rect 200662 633498 200746 633734
rect 200982 633498 236426 633734
rect 236662 633498 236746 633734
rect 236982 633498 272426 633734
rect 272662 633498 272746 633734
rect 272982 633498 308426 633734
rect 308662 633498 308746 633734
rect 308982 633498 344426 633734
rect 344662 633498 344746 633734
rect 344982 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 488426 633734
rect 488662 633498 488746 633734
rect 488982 633498 524426 633734
rect 524662 633498 524746 633734
rect 524982 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 592650 633734
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 52706 630334
rect 52942 630098 53026 630334
rect 53262 630098 88706 630334
rect 88942 630098 89026 630334
rect 89262 630098 124706 630334
rect 124942 630098 125026 630334
rect 125262 630098 160706 630334
rect 160942 630098 161026 630334
rect 161262 630098 196706 630334
rect 196942 630098 197026 630334
rect 197262 630098 232706 630334
rect 232942 630098 233026 630334
rect 233262 630098 268706 630334
rect 268942 630098 269026 630334
rect 269262 630098 304706 630334
rect 304942 630098 305026 630334
rect 305262 630098 340706 630334
rect 340942 630098 341026 630334
rect 341262 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 484706 630334
rect 484942 630098 485026 630334
rect 485262 630098 520706 630334
rect 520942 630098 521026 630334
rect 521262 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 592650 630334
rect -8726 630014 592650 630098
rect -8726 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 52706 630014
rect 52942 629778 53026 630014
rect 53262 629778 88706 630014
rect 88942 629778 89026 630014
rect 89262 629778 124706 630014
rect 124942 629778 125026 630014
rect 125262 629778 160706 630014
rect 160942 629778 161026 630014
rect 161262 629778 196706 630014
rect 196942 629778 197026 630014
rect 197262 629778 232706 630014
rect 232942 629778 233026 630014
rect 233262 629778 268706 630014
rect 268942 629778 269026 630014
rect 269262 629778 304706 630014
rect 304942 629778 305026 630014
rect 305262 629778 340706 630014
rect 340942 629778 341026 630014
rect 341262 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 484706 630014
rect 484942 629778 485026 630014
rect 485262 629778 520706 630014
rect 520942 629778 521026 630014
rect 521262 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 592650 630014
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 592650 626294
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 592650 622894
rect -8726 622574 592650 622658
rect -8726 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 592650 622574
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 592650 619174
rect -8726 618854 592650 618938
rect -8726 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 592650 618854
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 605494 592650 605526
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 63866 605494
rect 64102 605258 64186 605494
rect 64422 605258 99866 605494
rect 100102 605258 100186 605494
rect 100422 605258 135866 605494
rect 136102 605258 136186 605494
rect 136422 605258 171866 605494
rect 172102 605258 172186 605494
rect 172422 605258 207866 605494
rect 208102 605258 208186 605494
rect 208422 605258 243866 605494
rect 244102 605258 244186 605494
rect 244422 605258 279866 605494
rect 280102 605258 280186 605494
rect 280422 605258 315866 605494
rect 316102 605258 316186 605494
rect 316422 605258 351866 605494
rect 352102 605258 352186 605494
rect 352422 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 459866 605494
rect 460102 605258 460186 605494
rect 460422 605258 495866 605494
rect 496102 605258 496186 605494
rect 496422 605258 531866 605494
rect 532102 605258 532186 605494
rect 532422 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect -8726 605174 592650 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 63866 605174
rect 64102 604938 64186 605174
rect 64422 604938 99866 605174
rect 100102 604938 100186 605174
rect 100422 604938 135866 605174
rect 136102 604938 136186 605174
rect 136422 604938 171866 605174
rect 172102 604938 172186 605174
rect 172422 604938 207866 605174
rect 208102 604938 208186 605174
rect 208422 604938 243866 605174
rect 244102 604938 244186 605174
rect 244422 604938 279866 605174
rect 280102 604938 280186 605174
rect 280422 604938 315866 605174
rect 316102 604938 316186 605174
rect 316422 604938 351866 605174
rect 352102 604938 352186 605174
rect 352422 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 459866 605174
rect 460102 604938 460186 605174
rect 460422 604938 495866 605174
rect 496102 604938 496186 605174
rect 496422 604938 531866 605174
rect 532102 604938 532186 605174
rect 532422 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect -8726 604906 592650 604938
rect -8726 601774 592650 601806
rect -8726 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 24146 601774
rect 24382 601538 24466 601774
rect 24702 601538 60146 601774
rect 60382 601538 60466 601774
rect 60702 601538 96146 601774
rect 96382 601538 96466 601774
rect 96702 601538 132146 601774
rect 132382 601538 132466 601774
rect 132702 601538 168146 601774
rect 168382 601538 168466 601774
rect 168702 601538 204146 601774
rect 204382 601538 204466 601774
rect 204702 601538 240146 601774
rect 240382 601538 240466 601774
rect 240702 601538 276146 601774
rect 276382 601538 276466 601774
rect 276702 601538 312146 601774
rect 312382 601538 312466 601774
rect 312702 601538 348146 601774
rect 348382 601538 348466 601774
rect 348702 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 492146 601774
rect 492382 601538 492466 601774
rect 492702 601538 528146 601774
rect 528382 601538 528466 601774
rect 528702 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 592650 601774
rect -8726 601454 592650 601538
rect -8726 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 24146 601454
rect 24382 601218 24466 601454
rect 24702 601218 60146 601454
rect 60382 601218 60466 601454
rect 60702 601218 96146 601454
rect 96382 601218 96466 601454
rect 96702 601218 132146 601454
rect 132382 601218 132466 601454
rect 132702 601218 168146 601454
rect 168382 601218 168466 601454
rect 168702 601218 204146 601454
rect 204382 601218 204466 601454
rect 204702 601218 240146 601454
rect 240382 601218 240466 601454
rect 240702 601218 276146 601454
rect 276382 601218 276466 601454
rect 276702 601218 312146 601454
rect 312382 601218 312466 601454
rect 312702 601218 348146 601454
rect 348382 601218 348466 601454
rect 348702 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 492146 601454
rect 492382 601218 492466 601454
rect 492702 601218 528146 601454
rect 528382 601218 528466 601454
rect 528702 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 592650 601454
rect -8726 601186 592650 601218
rect -8726 598054 592650 598086
rect -8726 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 56426 598054
rect 56662 597818 56746 598054
rect 56982 597818 92426 598054
rect 92662 597818 92746 598054
rect 92982 597818 128426 598054
rect 128662 597818 128746 598054
rect 128982 597818 164426 598054
rect 164662 597818 164746 598054
rect 164982 597818 200426 598054
rect 200662 597818 200746 598054
rect 200982 597818 236426 598054
rect 236662 597818 236746 598054
rect 236982 597818 272426 598054
rect 272662 597818 272746 598054
rect 272982 597818 308426 598054
rect 308662 597818 308746 598054
rect 308982 597818 344426 598054
rect 344662 597818 344746 598054
rect 344982 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 592650 598054
rect -8726 597734 592650 597818
rect -8726 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 56426 597734
rect 56662 597498 56746 597734
rect 56982 597498 92426 597734
rect 92662 597498 92746 597734
rect 92982 597498 128426 597734
rect 128662 597498 128746 597734
rect 128982 597498 164426 597734
rect 164662 597498 164746 597734
rect 164982 597498 200426 597734
rect 200662 597498 200746 597734
rect 200982 597498 236426 597734
rect 236662 597498 236746 597734
rect 236982 597498 272426 597734
rect 272662 597498 272746 597734
rect 272982 597498 308426 597734
rect 308662 597498 308746 597734
rect 308982 597498 344426 597734
rect 344662 597498 344746 597734
rect 344982 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 592650 597734
rect -8726 597466 592650 597498
rect -8726 594334 592650 594366
rect -8726 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 52706 594334
rect 52942 594098 53026 594334
rect 53262 594098 88706 594334
rect 88942 594098 89026 594334
rect 89262 594098 124706 594334
rect 124942 594098 125026 594334
rect 125262 594098 160706 594334
rect 160942 594098 161026 594334
rect 161262 594098 196706 594334
rect 196942 594098 197026 594334
rect 197262 594098 232706 594334
rect 232942 594098 233026 594334
rect 233262 594098 268706 594334
rect 268942 594098 269026 594334
rect 269262 594098 304706 594334
rect 304942 594098 305026 594334
rect 305262 594098 340706 594334
rect 340942 594098 341026 594334
rect 341262 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 592650 594334
rect -8726 594014 592650 594098
rect -8726 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 52706 594014
rect 52942 593778 53026 594014
rect 53262 593778 88706 594014
rect 88942 593778 89026 594014
rect 89262 593778 124706 594014
rect 124942 593778 125026 594014
rect 125262 593778 160706 594014
rect 160942 593778 161026 594014
rect 161262 593778 196706 594014
rect 196942 593778 197026 594014
rect 197262 593778 232706 594014
rect 232942 593778 233026 594014
rect 233262 593778 268706 594014
rect 268942 593778 269026 594014
rect 269262 593778 304706 594014
rect 304942 593778 305026 594014
rect 305262 593778 340706 594014
rect 340942 593778 341026 594014
rect 341262 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 592650 594014
rect -8726 593746 592650 593778
rect -8726 590614 592650 590646
rect -8726 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 592650 590294
rect -8726 590026 592650 590058
rect -8726 586894 592650 586926
rect -8726 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 592650 586894
rect -8726 586574 592650 586658
rect -8726 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 592650 586574
rect -8726 586306 592650 586338
rect -8726 583174 592650 583206
rect -8726 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 592650 583174
rect -8726 582854 592650 582938
rect -8726 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 592650 582854
rect -8726 582586 592650 582618
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 569494 592650 569526
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 63866 569494
rect 64102 569258 64186 569494
rect 64422 569258 99866 569494
rect 100102 569258 100186 569494
rect 100422 569258 135866 569494
rect 136102 569258 136186 569494
rect 136422 569258 171866 569494
rect 172102 569258 172186 569494
rect 172422 569258 207866 569494
rect 208102 569258 208186 569494
rect 208422 569258 243866 569494
rect 244102 569258 244186 569494
rect 244422 569258 279866 569494
rect 280102 569258 280186 569494
rect 280422 569258 315866 569494
rect 316102 569258 316186 569494
rect 316422 569258 351866 569494
rect 352102 569258 352186 569494
rect 352422 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect -8726 569174 592650 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 63866 569174
rect 64102 568938 64186 569174
rect 64422 568938 99866 569174
rect 100102 568938 100186 569174
rect 100422 568938 135866 569174
rect 136102 568938 136186 569174
rect 136422 568938 171866 569174
rect 172102 568938 172186 569174
rect 172422 568938 207866 569174
rect 208102 568938 208186 569174
rect 208422 568938 243866 569174
rect 244102 568938 244186 569174
rect 244422 568938 279866 569174
rect 280102 568938 280186 569174
rect 280422 568938 315866 569174
rect 316102 568938 316186 569174
rect 316422 568938 351866 569174
rect 352102 568938 352186 569174
rect 352422 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect -8726 568906 592650 568938
rect -8726 565774 592650 565806
rect -8726 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 24146 565774
rect 24382 565538 24466 565774
rect 24702 565538 60146 565774
rect 60382 565538 60466 565774
rect 60702 565538 96146 565774
rect 96382 565538 96466 565774
rect 96702 565538 132146 565774
rect 132382 565538 132466 565774
rect 132702 565538 168146 565774
rect 168382 565538 168466 565774
rect 168702 565538 204146 565774
rect 204382 565538 204466 565774
rect 204702 565538 240146 565774
rect 240382 565538 240466 565774
rect 240702 565538 276146 565774
rect 276382 565538 276466 565774
rect 276702 565538 312146 565774
rect 312382 565538 312466 565774
rect 312702 565538 348146 565774
rect 348382 565538 348466 565774
rect 348702 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 420146 565774
rect 420382 565538 420466 565774
rect 420702 565538 456146 565774
rect 456382 565538 456466 565774
rect 456702 565538 492146 565774
rect 492382 565538 492466 565774
rect 492702 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 592650 565774
rect -8726 565454 592650 565538
rect -8726 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 24146 565454
rect 24382 565218 24466 565454
rect 24702 565218 60146 565454
rect 60382 565218 60466 565454
rect 60702 565218 96146 565454
rect 96382 565218 96466 565454
rect 96702 565218 132146 565454
rect 132382 565218 132466 565454
rect 132702 565218 168146 565454
rect 168382 565218 168466 565454
rect 168702 565218 204146 565454
rect 204382 565218 204466 565454
rect 204702 565218 240146 565454
rect 240382 565218 240466 565454
rect 240702 565218 276146 565454
rect 276382 565218 276466 565454
rect 276702 565218 312146 565454
rect 312382 565218 312466 565454
rect 312702 565218 348146 565454
rect 348382 565218 348466 565454
rect 348702 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 420146 565454
rect 420382 565218 420466 565454
rect 420702 565218 456146 565454
rect 456382 565218 456466 565454
rect 456702 565218 492146 565454
rect 492382 565218 492466 565454
rect 492702 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 592650 565454
rect -8726 565186 592650 565218
rect -8726 562054 592650 562086
rect -8726 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 56426 562054
rect 56662 561818 56746 562054
rect 56982 561818 92426 562054
rect 92662 561818 92746 562054
rect 92982 561818 128426 562054
rect 128662 561818 128746 562054
rect 128982 561818 164426 562054
rect 164662 561818 164746 562054
rect 164982 561818 200426 562054
rect 200662 561818 200746 562054
rect 200982 561818 236426 562054
rect 236662 561818 236746 562054
rect 236982 561818 272426 562054
rect 272662 561818 272746 562054
rect 272982 561818 308426 562054
rect 308662 561818 308746 562054
rect 308982 561818 344426 562054
rect 344662 561818 344746 562054
rect 344982 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 592650 562054
rect -8726 561734 592650 561818
rect -8726 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 56426 561734
rect 56662 561498 56746 561734
rect 56982 561498 92426 561734
rect 92662 561498 92746 561734
rect 92982 561498 128426 561734
rect 128662 561498 128746 561734
rect 128982 561498 164426 561734
rect 164662 561498 164746 561734
rect 164982 561498 200426 561734
rect 200662 561498 200746 561734
rect 200982 561498 236426 561734
rect 236662 561498 236746 561734
rect 236982 561498 272426 561734
rect 272662 561498 272746 561734
rect 272982 561498 308426 561734
rect 308662 561498 308746 561734
rect 308982 561498 344426 561734
rect 344662 561498 344746 561734
rect 344982 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 592650 561734
rect -8726 561466 592650 561498
rect -8726 558334 592650 558366
rect -8726 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 52706 558334
rect 52942 558098 53026 558334
rect 53262 558098 88706 558334
rect 88942 558098 89026 558334
rect 89262 558098 124706 558334
rect 124942 558098 125026 558334
rect 125262 558098 160706 558334
rect 160942 558098 161026 558334
rect 161262 558098 196706 558334
rect 196942 558098 197026 558334
rect 197262 558098 232706 558334
rect 232942 558098 233026 558334
rect 233262 558098 268706 558334
rect 268942 558098 269026 558334
rect 269262 558098 304706 558334
rect 304942 558098 305026 558334
rect 305262 558098 340706 558334
rect 340942 558098 341026 558334
rect 341262 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 592650 558334
rect -8726 558014 592650 558098
rect -8726 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 52706 558014
rect 52942 557778 53026 558014
rect 53262 557778 88706 558014
rect 88942 557778 89026 558014
rect 89262 557778 124706 558014
rect 124942 557778 125026 558014
rect 125262 557778 160706 558014
rect 160942 557778 161026 558014
rect 161262 557778 196706 558014
rect 196942 557778 197026 558014
rect 197262 557778 232706 558014
rect 232942 557778 233026 558014
rect 233262 557778 268706 558014
rect 268942 557778 269026 558014
rect 269262 557778 304706 558014
rect 304942 557778 305026 558014
rect 305262 557778 340706 558014
rect 340942 557778 341026 558014
rect 341262 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 592650 558014
rect -8726 557746 592650 557778
rect -8726 554614 592650 554646
rect -8726 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 592650 554294
rect -8726 554026 592650 554058
rect -8726 550894 592650 550926
rect -8726 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 592650 550894
rect -8726 550574 592650 550658
rect -8726 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 592650 550574
rect -8726 550306 592650 550338
rect -8726 547174 592650 547206
rect -8726 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 592650 547174
rect -8726 546854 592650 546938
rect -8726 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 592650 546854
rect -8726 546586 592650 546618
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 533494 592650 533526
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 63866 533494
rect 64102 533258 64186 533494
rect 64422 533258 99866 533494
rect 100102 533258 100186 533494
rect 100422 533258 135866 533494
rect 136102 533258 136186 533494
rect 136422 533258 171866 533494
rect 172102 533258 172186 533494
rect 172422 533258 207866 533494
rect 208102 533258 208186 533494
rect 208422 533258 243866 533494
rect 244102 533258 244186 533494
rect 244422 533258 279866 533494
rect 280102 533258 280186 533494
rect 280422 533258 315866 533494
rect 316102 533258 316186 533494
rect 316422 533258 351866 533494
rect 352102 533258 352186 533494
rect 352422 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect -8726 533174 592650 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 63866 533174
rect 64102 532938 64186 533174
rect 64422 532938 99866 533174
rect 100102 532938 100186 533174
rect 100422 532938 135866 533174
rect 136102 532938 136186 533174
rect 136422 532938 171866 533174
rect 172102 532938 172186 533174
rect 172422 532938 207866 533174
rect 208102 532938 208186 533174
rect 208422 532938 243866 533174
rect 244102 532938 244186 533174
rect 244422 532938 279866 533174
rect 280102 532938 280186 533174
rect 280422 532938 315866 533174
rect 316102 532938 316186 533174
rect 316422 532938 351866 533174
rect 352102 532938 352186 533174
rect 352422 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect -8726 532906 592650 532938
rect -8726 529774 592650 529806
rect -8726 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 24146 529774
rect 24382 529538 24466 529774
rect 24702 529538 60146 529774
rect 60382 529538 60466 529774
rect 60702 529538 96146 529774
rect 96382 529538 96466 529774
rect 96702 529538 132146 529774
rect 132382 529538 132466 529774
rect 132702 529538 168146 529774
rect 168382 529538 168466 529774
rect 168702 529538 204146 529774
rect 204382 529538 204466 529774
rect 204702 529538 240146 529774
rect 240382 529538 240466 529774
rect 240702 529538 276146 529774
rect 276382 529538 276466 529774
rect 276702 529538 312146 529774
rect 312382 529538 312466 529774
rect 312702 529538 348146 529774
rect 348382 529538 348466 529774
rect 348702 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 592650 529774
rect -8726 529454 592650 529538
rect -8726 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 24146 529454
rect 24382 529218 24466 529454
rect 24702 529218 60146 529454
rect 60382 529218 60466 529454
rect 60702 529218 96146 529454
rect 96382 529218 96466 529454
rect 96702 529218 132146 529454
rect 132382 529218 132466 529454
rect 132702 529218 168146 529454
rect 168382 529218 168466 529454
rect 168702 529218 204146 529454
rect 204382 529218 204466 529454
rect 204702 529218 240146 529454
rect 240382 529218 240466 529454
rect 240702 529218 276146 529454
rect 276382 529218 276466 529454
rect 276702 529218 312146 529454
rect 312382 529218 312466 529454
rect 312702 529218 348146 529454
rect 348382 529218 348466 529454
rect 348702 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 592650 529454
rect -8726 529186 592650 529218
rect -8726 526054 592650 526086
rect -8726 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 56426 526054
rect 56662 525818 56746 526054
rect 56982 525818 92426 526054
rect 92662 525818 92746 526054
rect 92982 525818 128426 526054
rect 128662 525818 128746 526054
rect 128982 525818 164426 526054
rect 164662 525818 164746 526054
rect 164982 525818 200426 526054
rect 200662 525818 200746 526054
rect 200982 525818 236426 526054
rect 236662 525818 236746 526054
rect 236982 525818 272426 526054
rect 272662 525818 272746 526054
rect 272982 525818 308426 526054
rect 308662 525818 308746 526054
rect 308982 525818 344426 526054
rect 344662 525818 344746 526054
rect 344982 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 592650 526054
rect -8726 525734 592650 525818
rect -8726 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 56426 525734
rect 56662 525498 56746 525734
rect 56982 525498 92426 525734
rect 92662 525498 92746 525734
rect 92982 525498 128426 525734
rect 128662 525498 128746 525734
rect 128982 525498 164426 525734
rect 164662 525498 164746 525734
rect 164982 525498 200426 525734
rect 200662 525498 200746 525734
rect 200982 525498 236426 525734
rect 236662 525498 236746 525734
rect 236982 525498 272426 525734
rect 272662 525498 272746 525734
rect 272982 525498 308426 525734
rect 308662 525498 308746 525734
rect 308982 525498 344426 525734
rect 344662 525498 344746 525734
rect 344982 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 592650 525734
rect -8726 525466 592650 525498
rect -8726 522334 592650 522366
rect -8726 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 52706 522334
rect 52942 522098 53026 522334
rect 53262 522098 88706 522334
rect 88942 522098 89026 522334
rect 89262 522098 124706 522334
rect 124942 522098 125026 522334
rect 125262 522098 160706 522334
rect 160942 522098 161026 522334
rect 161262 522098 196706 522334
rect 196942 522098 197026 522334
rect 197262 522098 232706 522334
rect 232942 522098 233026 522334
rect 233262 522098 268706 522334
rect 268942 522098 269026 522334
rect 269262 522098 304706 522334
rect 304942 522098 305026 522334
rect 305262 522098 340706 522334
rect 340942 522098 341026 522334
rect 341262 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 448706 522334
rect 448942 522098 449026 522334
rect 449262 522098 484706 522334
rect 484942 522098 485026 522334
rect 485262 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 592650 522334
rect -8726 522014 592650 522098
rect -8726 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 52706 522014
rect 52942 521778 53026 522014
rect 53262 521778 88706 522014
rect 88942 521778 89026 522014
rect 89262 521778 124706 522014
rect 124942 521778 125026 522014
rect 125262 521778 160706 522014
rect 160942 521778 161026 522014
rect 161262 521778 196706 522014
rect 196942 521778 197026 522014
rect 197262 521778 232706 522014
rect 232942 521778 233026 522014
rect 233262 521778 268706 522014
rect 268942 521778 269026 522014
rect 269262 521778 304706 522014
rect 304942 521778 305026 522014
rect 305262 521778 340706 522014
rect 340942 521778 341026 522014
rect 341262 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 448706 522014
rect 448942 521778 449026 522014
rect 449262 521778 484706 522014
rect 484942 521778 485026 522014
rect 485262 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 592650 522014
rect -8726 521746 592650 521778
rect -8726 518614 592650 518646
rect -8726 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 592650 518294
rect -8726 518026 592650 518058
rect -8726 514894 592650 514926
rect -8726 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 592650 514894
rect -8726 514574 592650 514658
rect -8726 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 592650 514574
rect -8726 514306 592650 514338
rect -8726 511174 592650 511206
rect -8726 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 592650 511174
rect -8726 510854 592650 510938
rect -8726 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 592650 510854
rect -8726 510586 592650 510618
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 497494 592650 497526
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 63866 497494
rect 64102 497258 64186 497494
rect 64422 497258 99866 497494
rect 100102 497258 100186 497494
rect 100422 497258 135866 497494
rect 136102 497258 136186 497494
rect 136422 497258 171866 497494
rect 172102 497258 172186 497494
rect 172422 497258 207866 497494
rect 208102 497258 208186 497494
rect 208422 497258 243866 497494
rect 244102 497258 244186 497494
rect 244422 497258 279866 497494
rect 280102 497258 280186 497494
rect 280422 497258 315866 497494
rect 316102 497258 316186 497494
rect 316422 497258 351866 497494
rect 352102 497258 352186 497494
rect 352422 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect -8726 497174 592650 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 63866 497174
rect 64102 496938 64186 497174
rect 64422 496938 99866 497174
rect 100102 496938 100186 497174
rect 100422 496938 135866 497174
rect 136102 496938 136186 497174
rect 136422 496938 171866 497174
rect 172102 496938 172186 497174
rect 172422 496938 207866 497174
rect 208102 496938 208186 497174
rect 208422 496938 243866 497174
rect 244102 496938 244186 497174
rect 244422 496938 279866 497174
rect 280102 496938 280186 497174
rect 280422 496938 315866 497174
rect 316102 496938 316186 497174
rect 316422 496938 351866 497174
rect 352102 496938 352186 497174
rect 352422 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect -8726 496906 592650 496938
rect -8726 493774 592650 493806
rect -8726 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 24146 493774
rect 24382 493538 24466 493774
rect 24702 493538 60146 493774
rect 60382 493538 60466 493774
rect 60702 493538 96146 493774
rect 96382 493538 96466 493774
rect 96702 493538 132146 493774
rect 132382 493538 132466 493774
rect 132702 493538 168146 493774
rect 168382 493538 168466 493774
rect 168702 493538 204146 493774
rect 204382 493538 204466 493774
rect 204702 493538 240146 493774
rect 240382 493538 240466 493774
rect 240702 493538 276146 493774
rect 276382 493538 276466 493774
rect 276702 493538 312146 493774
rect 312382 493538 312466 493774
rect 312702 493538 348146 493774
rect 348382 493538 348466 493774
rect 348702 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 420146 493774
rect 420382 493538 420466 493774
rect 420702 493538 456146 493774
rect 456382 493538 456466 493774
rect 456702 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 592650 493774
rect -8726 493454 592650 493538
rect -8726 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 24146 493454
rect 24382 493218 24466 493454
rect 24702 493218 60146 493454
rect 60382 493218 60466 493454
rect 60702 493218 96146 493454
rect 96382 493218 96466 493454
rect 96702 493218 132146 493454
rect 132382 493218 132466 493454
rect 132702 493218 168146 493454
rect 168382 493218 168466 493454
rect 168702 493218 204146 493454
rect 204382 493218 204466 493454
rect 204702 493218 240146 493454
rect 240382 493218 240466 493454
rect 240702 493218 276146 493454
rect 276382 493218 276466 493454
rect 276702 493218 312146 493454
rect 312382 493218 312466 493454
rect 312702 493218 348146 493454
rect 348382 493218 348466 493454
rect 348702 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 420146 493454
rect 420382 493218 420466 493454
rect 420702 493218 456146 493454
rect 456382 493218 456466 493454
rect 456702 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 592650 493454
rect -8726 493186 592650 493218
rect -8726 490054 592650 490086
rect -8726 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 56426 490054
rect 56662 489818 56746 490054
rect 56982 489818 92426 490054
rect 92662 489818 92746 490054
rect 92982 489818 128426 490054
rect 128662 489818 128746 490054
rect 128982 489818 164426 490054
rect 164662 489818 164746 490054
rect 164982 489818 200426 490054
rect 200662 489818 200746 490054
rect 200982 489818 236426 490054
rect 236662 489818 236746 490054
rect 236982 489818 272426 490054
rect 272662 489818 272746 490054
rect 272982 489818 308426 490054
rect 308662 489818 308746 490054
rect 308982 489818 344426 490054
rect 344662 489818 344746 490054
rect 344982 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 416426 490054
rect 416662 489818 416746 490054
rect 416982 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 592650 490054
rect -8726 489734 592650 489818
rect -8726 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 56426 489734
rect 56662 489498 56746 489734
rect 56982 489498 92426 489734
rect 92662 489498 92746 489734
rect 92982 489498 128426 489734
rect 128662 489498 128746 489734
rect 128982 489498 164426 489734
rect 164662 489498 164746 489734
rect 164982 489498 200426 489734
rect 200662 489498 200746 489734
rect 200982 489498 236426 489734
rect 236662 489498 236746 489734
rect 236982 489498 272426 489734
rect 272662 489498 272746 489734
rect 272982 489498 308426 489734
rect 308662 489498 308746 489734
rect 308982 489498 344426 489734
rect 344662 489498 344746 489734
rect 344982 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 416426 489734
rect 416662 489498 416746 489734
rect 416982 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 592650 489734
rect -8726 489466 592650 489498
rect -8726 486334 592650 486366
rect -8726 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 52706 486334
rect 52942 486098 53026 486334
rect 53262 486098 88706 486334
rect 88942 486098 89026 486334
rect 89262 486098 124706 486334
rect 124942 486098 125026 486334
rect 125262 486098 160706 486334
rect 160942 486098 161026 486334
rect 161262 486098 196706 486334
rect 196942 486098 197026 486334
rect 197262 486098 232706 486334
rect 232942 486098 233026 486334
rect 233262 486098 268706 486334
rect 268942 486098 269026 486334
rect 269262 486098 304706 486334
rect 304942 486098 305026 486334
rect 305262 486098 340706 486334
rect 340942 486098 341026 486334
rect 341262 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 412706 486334
rect 412942 486098 413026 486334
rect 413262 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 592650 486334
rect -8726 486014 592650 486098
rect -8726 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 52706 486014
rect 52942 485778 53026 486014
rect 53262 485778 88706 486014
rect 88942 485778 89026 486014
rect 89262 485778 124706 486014
rect 124942 485778 125026 486014
rect 125262 485778 160706 486014
rect 160942 485778 161026 486014
rect 161262 485778 196706 486014
rect 196942 485778 197026 486014
rect 197262 485778 232706 486014
rect 232942 485778 233026 486014
rect 233262 485778 268706 486014
rect 268942 485778 269026 486014
rect 269262 485778 304706 486014
rect 304942 485778 305026 486014
rect 305262 485778 340706 486014
rect 340942 485778 341026 486014
rect 341262 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 412706 486014
rect 412942 485778 413026 486014
rect 413262 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 592650 486014
rect -8726 485746 592650 485778
rect -8726 482614 592650 482646
rect -8726 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 592650 482294
rect -8726 482026 592650 482058
rect -8726 478894 592650 478926
rect -8726 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 592650 478894
rect -8726 478574 592650 478658
rect -8726 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 592650 478574
rect -8726 478306 592650 478338
rect -8726 475174 592650 475206
rect -8726 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 592650 475174
rect -8726 474854 592650 474938
rect -8726 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 592650 474854
rect -8726 474586 592650 474618
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 461494 592650 461526
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 63866 461494
rect 64102 461258 64186 461494
rect 64422 461258 99866 461494
rect 100102 461258 100186 461494
rect 100422 461258 135866 461494
rect 136102 461258 136186 461494
rect 136422 461258 171866 461494
rect 172102 461258 172186 461494
rect 172422 461258 207866 461494
rect 208102 461258 208186 461494
rect 208422 461258 243866 461494
rect 244102 461258 244186 461494
rect 244422 461258 279866 461494
rect 280102 461258 280186 461494
rect 280422 461258 315866 461494
rect 316102 461258 316186 461494
rect 316422 461258 351866 461494
rect 352102 461258 352186 461494
rect 352422 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect -8726 461174 592650 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 63866 461174
rect 64102 460938 64186 461174
rect 64422 460938 99866 461174
rect 100102 460938 100186 461174
rect 100422 460938 135866 461174
rect 136102 460938 136186 461174
rect 136422 460938 171866 461174
rect 172102 460938 172186 461174
rect 172422 460938 207866 461174
rect 208102 460938 208186 461174
rect 208422 460938 243866 461174
rect 244102 460938 244186 461174
rect 244422 460938 279866 461174
rect 280102 460938 280186 461174
rect 280422 460938 315866 461174
rect 316102 460938 316186 461174
rect 316422 460938 351866 461174
rect 352102 460938 352186 461174
rect 352422 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect -8726 460906 592650 460938
rect -8726 457774 592650 457806
rect -8726 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 24146 457774
rect 24382 457538 24466 457774
rect 24702 457538 60146 457774
rect 60382 457538 60466 457774
rect 60702 457538 96146 457774
rect 96382 457538 96466 457774
rect 96702 457538 132146 457774
rect 132382 457538 132466 457774
rect 132702 457538 168146 457774
rect 168382 457538 168466 457774
rect 168702 457538 204146 457774
rect 204382 457538 204466 457774
rect 204702 457538 240146 457774
rect 240382 457538 240466 457774
rect 240702 457538 276146 457774
rect 276382 457538 276466 457774
rect 276702 457538 312146 457774
rect 312382 457538 312466 457774
rect 312702 457538 348146 457774
rect 348382 457538 348466 457774
rect 348702 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 420146 457774
rect 420382 457538 420466 457774
rect 420702 457538 456146 457774
rect 456382 457538 456466 457774
rect 456702 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 592650 457774
rect -8726 457454 592650 457538
rect -8726 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 24146 457454
rect 24382 457218 24466 457454
rect 24702 457218 60146 457454
rect 60382 457218 60466 457454
rect 60702 457218 96146 457454
rect 96382 457218 96466 457454
rect 96702 457218 132146 457454
rect 132382 457218 132466 457454
rect 132702 457218 168146 457454
rect 168382 457218 168466 457454
rect 168702 457218 204146 457454
rect 204382 457218 204466 457454
rect 204702 457218 240146 457454
rect 240382 457218 240466 457454
rect 240702 457218 276146 457454
rect 276382 457218 276466 457454
rect 276702 457218 312146 457454
rect 312382 457218 312466 457454
rect 312702 457218 348146 457454
rect 348382 457218 348466 457454
rect 348702 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 420146 457454
rect 420382 457218 420466 457454
rect 420702 457218 456146 457454
rect 456382 457218 456466 457454
rect 456702 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 592650 457454
rect -8726 457186 592650 457218
rect -8726 454054 592650 454086
rect -8726 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 56426 454054
rect 56662 453818 56746 454054
rect 56982 453818 92426 454054
rect 92662 453818 92746 454054
rect 92982 453818 128426 454054
rect 128662 453818 128746 454054
rect 128982 453818 164426 454054
rect 164662 453818 164746 454054
rect 164982 453818 200426 454054
rect 200662 453818 200746 454054
rect 200982 453818 236426 454054
rect 236662 453818 236746 454054
rect 236982 453818 272426 454054
rect 272662 453818 272746 454054
rect 272982 453818 308426 454054
rect 308662 453818 308746 454054
rect 308982 453818 344426 454054
rect 344662 453818 344746 454054
rect 344982 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 416426 454054
rect 416662 453818 416746 454054
rect 416982 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 453818 488426 454054
rect 488662 453818 488746 454054
rect 488982 453818 524426 454054
rect 524662 453818 524746 454054
rect 524982 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 592650 454054
rect -8726 453734 592650 453818
rect -8726 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 56426 453734
rect 56662 453498 56746 453734
rect 56982 453498 92426 453734
rect 92662 453498 92746 453734
rect 92982 453498 128426 453734
rect 128662 453498 128746 453734
rect 128982 453498 164426 453734
rect 164662 453498 164746 453734
rect 164982 453498 200426 453734
rect 200662 453498 200746 453734
rect 200982 453498 236426 453734
rect 236662 453498 236746 453734
rect 236982 453498 272426 453734
rect 272662 453498 272746 453734
rect 272982 453498 308426 453734
rect 308662 453498 308746 453734
rect 308982 453498 344426 453734
rect 344662 453498 344746 453734
rect 344982 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 416426 453734
rect 416662 453498 416746 453734
rect 416982 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 488426 453734
rect 488662 453498 488746 453734
rect 488982 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 592650 453734
rect -8726 453466 592650 453498
rect -8726 450334 592650 450366
rect -8726 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 52706 450334
rect 52942 450098 53026 450334
rect 53262 450098 88706 450334
rect 88942 450098 89026 450334
rect 89262 450098 124706 450334
rect 124942 450098 125026 450334
rect 125262 450098 160706 450334
rect 160942 450098 161026 450334
rect 161262 450098 196706 450334
rect 196942 450098 197026 450334
rect 197262 450098 232706 450334
rect 232942 450098 233026 450334
rect 233262 450098 268706 450334
rect 268942 450098 269026 450334
rect 269262 450098 304706 450334
rect 304942 450098 305026 450334
rect 305262 450098 340706 450334
rect 340942 450098 341026 450334
rect 341262 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 412706 450334
rect 412942 450098 413026 450334
rect 413262 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 592650 450334
rect -8726 450014 592650 450098
rect -8726 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 52706 450014
rect 52942 449778 53026 450014
rect 53262 449778 88706 450014
rect 88942 449778 89026 450014
rect 89262 449778 124706 450014
rect 124942 449778 125026 450014
rect 125262 449778 160706 450014
rect 160942 449778 161026 450014
rect 161262 449778 196706 450014
rect 196942 449778 197026 450014
rect 197262 449778 232706 450014
rect 232942 449778 233026 450014
rect 233262 449778 268706 450014
rect 268942 449778 269026 450014
rect 269262 449778 304706 450014
rect 304942 449778 305026 450014
rect 305262 449778 340706 450014
rect 340942 449778 341026 450014
rect 341262 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 412706 450014
rect 412942 449778 413026 450014
rect 413262 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 592650 450014
rect -8726 449746 592650 449778
rect -8726 446614 592650 446646
rect -8726 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 592650 446294
rect -8726 446026 592650 446058
rect -8726 442894 592650 442926
rect -8726 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 592650 442894
rect -8726 442574 592650 442658
rect -8726 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 592650 442574
rect -8726 442306 592650 442338
rect -8726 439174 592650 439206
rect -8726 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 592650 439174
rect -8726 438854 592650 438938
rect -8726 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 592650 438854
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 425494 592650 425526
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 63866 425494
rect 64102 425258 64186 425494
rect 64422 425258 99866 425494
rect 100102 425258 100186 425494
rect 100422 425258 135866 425494
rect 136102 425258 136186 425494
rect 136422 425258 171866 425494
rect 172102 425258 172186 425494
rect 172422 425258 207866 425494
rect 208102 425258 208186 425494
rect 208422 425258 243866 425494
rect 244102 425258 244186 425494
rect 244422 425258 279866 425494
rect 280102 425258 280186 425494
rect 280422 425258 315866 425494
rect 316102 425258 316186 425494
rect 316422 425258 351866 425494
rect 352102 425258 352186 425494
rect 352422 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 423866 425494
rect 424102 425258 424186 425494
rect 424422 425258 459866 425494
rect 460102 425258 460186 425494
rect 460422 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect -8726 425174 592650 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 63866 425174
rect 64102 424938 64186 425174
rect 64422 424938 99866 425174
rect 100102 424938 100186 425174
rect 100422 424938 135866 425174
rect 136102 424938 136186 425174
rect 136422 424938 171866 425174
rect 172102 424938 172186 425174
rect 172422 424938 207866 425174
rect 208102 424938 208186 425174
rect 208422 424938 243866 425174
rect 244102 424938 244186 425174
rect 244422 424938 279866 425174
rect 280102 424938 280186 425174
rect 280422 424938 315866 425174
rect 316102 424938 316186 425174
rect 316422 424938 351866 425174
rect 352102 424938 352186 425174
rect 352422 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 423866 425174
rect 424102 424938 424186 425174
rect 424422 424938 459866 425174
rect 460102 424938 460186 425174
rect 460422 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect -8726 424906 592650 424938
rect -8726 421774 592650 421806
rect -8726 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 24146 421774
rect 24382 421538 24466 421774
rect 24702 421538 60146 421774
rect 60382 421538 60466 421774
rect 60702 421538 96146 421774
rect 96382 421538 96466 421774
rect 96702 421538 132146 421774
rect 132382 421538 132466 421774
rect 132702 421538 168146 421774
rect 168382 421538 168466 421774
rect 168702 421538 204146 421774
rect 204382 421538 204466 421774
rect 204702 421538 240146 421774
rect 240382 421538 240466 421774
rect 240702 421538 276146 421774
rect 276382 421538 276466 421774
rect 276702 421538 312146 421774
rect 312382 421538 312466 421774
rect 312702 421538 348146 421774
rect 348382 421538 348466 421774
rect 348702 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 420146 421774
rect 420382 421538 420466 421774
rect 420702 421538 456146 421774
rect 456382 421538 456466 421774
rect 456702 421538 492146 421774
rect 492382 421538 492466 421774
rect 492702 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 592650 421774
rect -8726 421454 592650 421538
rect -8726 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 24146 421454
rect 24382 421218 24466 421454
rect 24702 421218 60146 421454
rect 60382 421218 60466 421454
rect 60702 421218 96146 421454
rect 96382 421218 96466 421454
rect 96702 421218 132146 421454
rect 132382 421218 132466 421454
rect 132702 421218 168146 421454
rect 168382 421218 168466 421454
rect 168702 421218 204146 421454
rect 204382 421218 204466 421454
rect 204702 421218 240146 421454
rect 240382 421218 240466 421454
rect 240702 421218 276146 421454
rect 276382 421218 276466 421454
rect 276702 421218 312146 421454
rect 312382 421218 312466 421454
rect 312702 421218 348146 421454
rect 348382 421218 348466 421454
rect 348702 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 420146 421454
rect 420382 421218 420466 421454
rect 420702 421218 456146 421454
rect 456382 421218 456466 421454
rect 456702 421218 492146 421454
rect 492382 421218 492466 421454
rect 492702 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 592650 421454
rect -8726 421186 592650 421218
rect -8726 418054 592650 418086
rect -8726 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 56426 418054
rect 56662 417818 56746 418054
rect 56982 417818 92426 418054
rect 92662 417818 92746 418054
rect 92982 417818 128426 418054
rect 128662 417818 128746 418054
rect 128982 417818 164426 418054
rect 164662 417818 164746 418054
rect 164982 417818 200426 418054
rect 200662 417818 200746 418054
rect 200982 417818 236426 418054
rect 236662 417818 236746 418054
rect 236982 417818 272426 418054
rect 272662 417818 272746 418054
rect 272982 417818 308426 418054
rect 308662 417818 308746 418054
rect 308982 417818 344426 418054
rect 344662 417818 344746 418054
rect 344982 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 416426 418054
rect 416662 417818 416746 418054
rect 416982 417818 452426 418054
rect 452662 417818 452746 418054
rect 452982 417818 488426 418054
rect 488662 417818 488746 418054
rect 488982 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 592650 418054
rect -8726 417734 592650 417818
rect -8726 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 56426 417734
rect 56662 417498 56746 417734
rect 56982 417498 92426 417734
rect 92662 417498 92746 417734
rect 92982 417498 128426 417734
rect 128662 417498 128746 417734
rect 128982 417498 164426 417734
rect 164662 417498 164746 417734
rect 164982 417498 200426 417734
rect 200662 417498 200746 417734
rect 200982 417498 236426 417734
rect 236662 417498 236746 417734
rect 236982 417498 272426 417734
rect 272662 417498 272746 417734
rect 272982 417498 308426 417734
rect 308662 417498 308746 417734
rect 308982 417498 344426 417734
rect 344662 417498 344746 417734
rect 344982 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 416426 417734
rect 416662 417498 416746 417734
rect 416982 417498 452426 417734
rect 452662 417498 452746 417734
rect 452982 417498 488426 417734
rect 488662 417498 488746 417734
rect 488982 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 592650 417734
rect -8726 417466 592650 417498
rect -8726 414334 592650 414366
rect -8726 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 52706 414334
rect 52942 414098 53026 414334
rect 53262 414098 88706 414334
rect 88942 414098 89026 414334
rect 89262 414098 124706 414334
rect 124942 414098 125026 414334
rect 125262 414098 160706 414334
rect 160942 414098 161026 414334
rect 161262 414098 196706 414334
rect 196942 414098 197026 414334
rect 197262 414098 232706 414334
rect 232942 414098 233026 414334
rect 233262 414098 268706 414334
rect 268942 414098 269026 414334
rect 269262 414098 304706 414334
rect 304942 414098 305026 414334
rect 305262 414098 340706 414334
rect 340942 414098 341026 414334
rect 341262 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 412706 414334
rect 412942 414098 413026 414334
rect 413262 414098 448706 414334
rect 448942 414098 449026 414334
rect 449262 414098 484706 414334
rect 484942 414098 485026 414334
rect 485262 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 592650 414334
rect -8726 414014 592650 414098
rect -8726 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 52706 414014
rect 52942 413778 53026 414014
rect 53262 413778 88706 414014
rect 88942 413778 89026 414014
rect 89262 413778 124706 414014
rect 124942 413778 125026 414014
rect 125262 413778 160706 414014
rect 160942 413778 161026 414014
rect 161262 413778 196706 414014
rect 196942 413778 197026 414014
rect 197262 413778 232706 414014
rect 232942 413778 233026 414014
rect 233262 413778 268706 414014
rect 268942 413778 269026 414014
rect 269262 413778 304706 414014
rect 304942 413778 305026 414014
rect 305262 413778 340706 414014
rect 340942 413778 341026 414014
rect 341262 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 412706 414014
rect 412942 413778 413026 414014
rect 413262 413778 448706 414014
rect 448942 413778 449026 414014
rect 449262 413778 484706 414014
rect 484942 413778 485026 414014
rect 485262 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 592650 414014
rect -8726 413746 592650 413778
rect -8726 410614 592650 410646
rect -8726 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 592650 410294
rect -8726 410026 592650 410058
rect -8726 406894 592650 406926
rect -8726 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 592650 406894
rect -8726 406574 592650 406658
rect -8726 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 592650 406574
rect -8726 406306 592650 406338
rect -8726 403174 592650 403206
rect -8726 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 592650 403174
rect -8726 402854 592650 402938
rect -8726 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 592650 402854
rect -8726 402586 592650 402618
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 389494 592650 389526
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 63866 389494
rect 64102 389258 64186 389494
rect 64422 389258 99866 389494
rect 100102 389258 100186 389494
rect 100422 389258 135866 389494
rect 136102 389258 136186 389494
rect 136422 389258 171866 389494
rect 172102 389258 172186 389494
rect 172422 389258 207866 389494
rect 208102 389258 208186 389494
rect 208422 389258 243866 389494
rect 244102 389258 244186 389494
rect 244422 389258 279866 389494
rect 280102 389258 280186 389494
rect 280422 389258 315866 389494
rect 316102 389258 316186 389494
rect 316422 389258 351866 389494
rect 352102 389258 352186 389494
rect 352422 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 423866 389494
rect 424102 389258 424186 389494
rect 424422 389258 459866 389494
rect 460102 389258 460186 389494
rect 460422 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect -8726 389174 592650 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 63866 389174
rect 64102 388938 64186 389174
rect 64422 388938 99866 389174
rect 100102 388938 100186 389174
rect 100422 388938 135866 389174
rect 136102 388938 136186 389174
rect 136422 388938 171866 389174
rect 172102 388938 172186 389174
rect 172422 388938 207866 389174
rect 208102 388938 208186 389174
rect 208422 388938 243866 389174
rect 244102 388938 244186 389174
rect 244422 388938 279866 389174
rect 280102 388938 280186 389174
rect 280422 388938 315866 389174
rect 316102 388938 316186 389174
rect 316422 388938 351866 389174
rect 352102 388938 352186 389174
rect 352422 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 423866 389174
rect 424102 388938 424186 389174
rect 424422 388938 459866 389174
rect 460102 388938 460186 389174
rect 460422 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect -8726 388906 592650 388938
rect -8726 385774 592650 385806
rect -8726 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 24146 385774
rect 24382 385538 24466 385774
rect 24702 385538 60146 385774
rect 60382 385538 60466 385774
rect 60702 385538 96146 385774
rect 96382 385538 96466 385774
rect 96702 385538 132146 385774
rect 132382 385538 132466 385774
rect 132702 385538 168146 385774
rect 168382 385538 168466 385774
rect 168702 385538 204146 385774
rect 204382 385538 204466 385774
rect 204702 385538 240146 385774
rect 240382 385538 240466 385774
rect 240702 385538 276146 385774
rect 276382 385538 276466 385774
rect 276702 385538 312146 385774
rect 312382 385538 312466 385774
rect 312702 385538 348146 385774
rect 348382 385538 348466 385774
rect 348702 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 492146 385774
rect 492382 385538 492466 385774
rect 492702 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 592650 385774
rect -8726 385454 592650 385538
rect -8726 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 24146 385454
rect 24382 385218 24466 385454
rect 24702 385218 60146 385454
rect 60382 385218 60466 385454
rect 60702 385218 96146 385454
rect 96382 385218 96466 385454
rect 96702 385218 132146 385454
rect 132382 385218 132466 385454
rect 132702 385218 168146 385454
rect 168382 385218 168466 385454
rect 168702 385218 204146 385454
rect 204382 385218 204466 385454
rect 204702 385218 240146 385454
rect 240382 385218 240466 385454
rect 240702 385218 276146 385454
rect 276382 385218 276466 385454
rect 276702 385218 312146 385454
rect 312382 385218 312466 385454
rect 312702 385218 348146 385454
rect 348382 385218 348466 385454
rect 348702 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 492146 385454
rect 492382 385218 492466 385454
rect 492702 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 592650 385454
rect -8726 385186 592650 385218
rect -8726 382054 592650 382086
rect -8726 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 56426 382054
rect 56662 381818 56746 382054
rect 56982 381818 92426 382054
rect 92662 381818 92746 382054
rect 92982 381818 128426 382054
rect 128662 381818 128746 382054
rect 128982 381818 164426 382054
rect 164662 381818 164746 382054
rect 164982 381818 200426 382054
rect 200662 381818 200746 382054
rect 200982 381818 236426 382054
rect 236662 381818 236746 382054
rect 236982 381818 272426 382054
rect 272662 381818 272746 382054
rect 272982 381818 308426 382054
rect 308662 381818 308746 382054
rect 308982 381818 344426 382054
rect 344662 381818 344746 382054
rect 344982 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 488426 382054
rect 488662 381818 488746 382054
rect 488982 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 592650 382054
rect -8726 381734 592650 381818
rect -8726 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 56426 381734
rect 56662 381498 56746 381734
rect 56982 381498 92426 381734
rect 92662 381498 92746 381734
rect 92982 381498 128426 381734
rect 128662 381498 128746 381734
rect 128982 381498 164426 381734
rect 164662 381498 164746 381734
rect 164982 381498 200426 381734
rect 200662 381498 200746 381734
rect 200982 381498 236426 381734
rect 236662 381498 236746 381734
rect 236982 381498 272426 381734
rect 272662 381498 272746 381734
rect 272982 381498 308426 381734
rect 308662 381498 308746 381734
rect 308982 381498 344426 381734
rect 344662 381498 344746 381734
rect 344982 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 488426 381734
rect 488662 381498 488746 381734
rect 488982 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 592650 381734
rect -8726 381466 592650 381498
rect -8726 378334 592650 378366
rect -8726 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 52706 378334
rect 52942 378098 53026 378334
rect 53262 378098 88706 378334
rect 88942 378098 89026 378334
rect 89262 378098 124706 378334
rect 124942 378098 125026 378334
rect 125262 378098 160706 378334
rect 160942 378098 161026 378334
rect 161262 378098 196706 378334
rect 196942 378098 197026 378334
rect 197262 378098 232706 378334
rect 232942 378098 233026 378334
rect 233262 378098 268706 378334
rect 268942 378098 269026 378334
rect 269262 378098 304706 378334
rect 304942 378098 305026 378334
rect 305262 378098 340706 378334
rect 340942 378098 341026 378334
rect 341262 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 484706 378334
rect 484942 378098 485026 378334
rect 485262 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378098 556706 378334
rect 556942 378098 557026 378334
rect 557262 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 592650 378334
rect -8726 378014 592650 378098
rect -8726 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 52706 378014
rect 52942 377778 53026 378014
rect 53262 377778 88706 378014
rect 88942 377778 89026 378014
rect 89262 377778 124706 378014
rect 124942 377778 125026 378014
rect 125262 377778 160706 378014
rect 160942 377778 161026 378014
rect 161262 377778 196706 378014
rect 196942 377778 197026 378014
rect 197262 377778 232706 378014
rect 232942 377778 233026 378014
rect 233262 377778 268706 378014
rect 268942 377778 269026 378014
rect 269262 377778 304706 378014
rect 304942 377778 305026 378014
rect 305262 377778 340706 378014
rect 340942 377778 341026 378014
rect 341262 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 484706 378014
rect 484942 377778 485026 378014
rect 485262 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 377778 556706 378014
rect 556942 377778 557026 378014
rect 557262 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 592650 378014
rect -8726 377746 592650 377778
rect -8726 374614 592650 374646
rect -8726 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 592650 374294
rect -8726 374026 592650 374058
rect -8726 370894 592650 370926
rect -8726 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 592650 370894
rect -8726 370574 592650 370658
rect -8726 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 592650 370574
rect -8726 370306 592650 370338
rect -8726 367174 592650 367206
rect -8726 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 592650 367174
rect -8726 366854 592650 366938
rect -8726 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 592650 366854
rect -8726 366586 592650 366618
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 353494 592650 353526
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 63866 353494
rect 64102 353258 64186 353494
rect 64422 353258 99866 353494
rect 100102 353258 100186 353494
rect 100422 353258 135866 353494
rect 136102 353258 136186 353494
rect 136422 353258 171866 353494
rect 172102 353258 172186 353494
rect 172422 353258 207866 353494
rect 208102 353258 208186 353494
rect 208422 353258 243866 353494
rect 244102 353258 244186 353494
rect 244422 353258 279866 353494
rect 280102 353258 280186 353494
rect 280422 353258 315866 353494
rect 316102 353258 316186 353494
rect 316422 353258 351866 353494
rect 352102 353258 352186 353494
rect 352422 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 495866 353494
rect 496102 353258 496186 353494
rect 496422 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect -8726 353174 592650 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 63866 353174
rect 64102 352938 64186 353174
rect 64422 352938 99866 353174
rect 100102 352938 100186 353174
rect 100422 352938 135866 353174
rect 136102 352938 136186 353174
rect 136422 352938 171866 353174
rect 172102 352938 172186 353174
rect 172422 352938 207866 353174
rect 208102 352938 208186 353174
rect 208422 352938 243866 353174
rect 244102 352938 244186 353174
rect 244422 352938 279866 353174
rect 280102 352938 280186 353174
rect 280422 352938 315866 353174
rect 316102 352938 316186 353174
rect 316422 352938 351866 353174
rect 352102 352938 352186 353174
rect 352422 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 495866 353174
rect 496102 352938 496186 353174
rect 496422 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect -8726 352906 592650 352938
rect -8726 349774 592650 349806
rect -8726 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 24146 349774
rect 24382 349538 24466 349774
rect 24702 349538 60146 349774
rect 60382 349538 60466 349774
rect 60702 349538 96146 349774
rect 96382 349538 96466 349774
rect 96702 349538 132146 349774
rect 132382 349538 132466 349774
rect 132702 349538 168146 349774
rect 168382 349538 168466 349774
rect 168702 349538 204146 349774
rect 204382 349538 204466 349774
rect 204702 349538 240146 349774
rect 240382 349538 240466 349774
rect 240702 349538 276146 349774
rect 276382 349538 276466 349774
rect 276702 349538 312146 349774
rect 312382 349538 312466 349774
rect 312702 349538 348146 349774
rect 348382 349538 348466 349774
rect 348702 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 492146 349774
rect 492382 349538 492466 349774
rect 492702 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 592650 349774
rect -8726 349454 592650 349538
rect -8726 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 24146 349454
rect 24382 349218 24466 349454
rect 24702 349218 60146 349454
rect 60382 349218 60466 349454
rect 60702 349218 96146 349454
rect 96382 349218 96466 349454
rect 96702 349218 132146 349454
rect 132382 349218 132466 349454
rect 132702 349218 168146 349454
rect 168382 349218 168466 349454
rect 168702 349218 204146 349454
rect 204382 349218 204466 349454
rect 204702 349218 240146 349454
rect 240382 349218 240466 349454
rect 240702 349218 276146 349454
rect 276382 349218 276466 349454
rect 276702 349218 312146 349454
rect 312382 349218 312466 349454
rect 312702 349218 348146 349454
rect 348382 349218 348466 349454
rect 348702 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 492146 349454
rect 492382 349218 492466 349454
rect 492702 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 592650 349454
rect -8726 349186 592650 349218
rect -8726 346054 592650 346086
rect -8726 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 56426 346054
rect 56662 345818 56746 346054
rect 56982 345818 92426 346054
rect 92662 345818 92746 346054
rect 92982 345818 128426 346054
rect 128662 345818 128746 346054
rect 128982 345818 164426 346054
rect 164662 345818 164746 346054
rect 164982 345818 200426 346054
rect 200662 345818 200746 346054
rect 200982 345818 236426 346054
rect 236662 345818 236746 346054
rect 236982 345818 272426 346054
rect 272662 345818 272746 346054
rect 272982 345818 308426 346054
rect 308662 345818 308746 346054
rect 308982 345818 344426 346054
rect 344662 345818 344746 346054
rect 344982 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 488426 346054
rect 488662 345818 488746 346054
rect 488982 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 592650 346054
rect -8726 345734 592650 345818
rect -8726 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 56426 345734
rect 56662 345498 56746 345734
rect 56982 345498 92426 345734
rect 92662 345498 92746 345734
rect 92982 345498 128426 345734
rect 128662 345498 128746 345734
rect 128982 345498 164426 345734
rect 164662 345498 164746 345734
rect 164982 345498 200426 345734
rect 200662 345498 200746 345734
rect 200982 345498 236426 345734
rect 236662 345498 236746 345734
rect 236982 345498 272426 345734
rect 272662 345498 272746 345734
rect 272982 345498 308426 345734
rect 308662 345498 308746 345734
rect 308982 345498 344426 345734
rect 344662 345498 344746 345734
rect 344982 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 488426 345734
rect 488662 345498 488746 345734
rect 488982 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 592650 345734
rect -8726 345466 592650 345498
rect -8726 342334 592650 342366
rect -8726 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 52706 342334
rect 52942 342098 53026 342334
rect 53262 342098 88706 342334
rect 88942 342098 89026 342334
rect 89262 342098 124706 342334
rect 124942 342098 125026 342334
rect 125262 342098 160706 342334
rect 160942 342098 161026 342334
rect 161262 342098 196706 342334
rect 196942 342098 197026 342334
rect 197262 342098 232706 342334
rect 232942 342098 233026 342334
rect 233262 342098 268706 342334
rect 268942 342098 269026 342334
rect 269262 342098 304706 342334
rect 304942 342098 305026 342334
rect 305262 342098 340706 342334
rect 340942 342098 341026 342334
rect 341262 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 484706 342334
rect 484942 342098 485026 342334
rect 485262 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 592650 342334
rect -8726 342014 592650 342098
rect -8726 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 52706 342014
rect 52942 341778 53026 342014
rect 53262 341778 88706 342014
rect 88942 341778 89026 342014
rect 89262 341778 124706 342014
rect 124942 341778 125026 342014
rect 125262 341778 160706 342014
rect 160942 341778 161026 342014
rect 161262 341778 196706 342014
rect 196942 341778 197026 342014
rect 197262 341778 232706 342014
rect 232942 341778 233026 342014
rect 233262 341778 268706 342014
rect 268942 341778 269026 342014
rect 269262 341778 304706 342014
rect 304942 341778 305026 342014
rect 305262 341778 340706 342014
rect 340942 341778 341026 342014
rect 341262 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 484706 342014
rect 484942 341778 485026 342014
rect 485262 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 592650 342014
rect -8726 341746 592650 341778
rect -8726 338614 592650 338646
rect -8726 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 592650 338294
rect -8726 338026 592650 338058
rect -8726 334894 592650 334926
rect -8726 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 592650 334894
rect -8726 334574 592650 334658
rect -8726 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 592650 334574
rect -8726 334306 592650 334338
rect -8726 331174 592650 331206
rect -8726 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 592650 331174
rect -8726 330854 592650 330938
rect -8726 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 592650 330854
rect -8726 330586 592650 330618
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 317494 592650 317526
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 63866 317494
rect 64102 317258 64186 317494
rect 64422 317258 99866 317494
rect 100102 317258 100186 317494
rect 100422 317258 135866 317494
rect 136102 317258 136186 317494
rect 136422 317258 171866 317494
rect 172102 317258 172186 317494
rect 172422 317258 207866 317494
rect 208102 317258 208186 317494
rect 208422 317258 243866 317494
rect 244102 317258 244186 317494
rect 244422 317258 279866 317494
rect 280102 317258 280186 317494
rect 280422 317258 315866 317494
rect 316102 317258 316186 317494
rect 316422 317258 351866 317494
rect 352102 317258 352186 317494
rect 352422 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect -8726 317174 592650 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 63866 317174
rect 64102 316938 64186 317174
rect 64422 316938 99866 317174
rect 100102 316938 100186 317174
rect 100422 316938 135866 317174
rect 136102 316938 136186 317174
rect 136422 316938 171866 317174
rect 172102 316938 172186 317174
rect 172422 316938 207866 317174
rect 208102 316938 208186 317174
rect 208422 316938 243866 317174
rect 244102 316938 244186 317174
rect 244422 316938 279866 317174
rect 280102 316938 280186 317174
rect 280422 316938 315866 317174
rect 316102 316938 316186 317174
rect 316422 316938 351866 317174
rect 352102 316938 352186 317174
rect 352422 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect -8726 316906 592650 316938
rect -8726 313774 592650 313806
rect -8726 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 24146 313774
rect 24382 313538 24466 313774
rect 24702 313538 60146 313774
rect 60382 313538 60466 313774
rect 60702 313538 96146 313774
rect 96382 313538 96466 313774
rect 96702 313538 132146 313774
rect 132382 313538 132466 313774
rect 132702 313538 168146 313774
rect 168382 313538 168466 313774
rect 168702 313538 204146 313774
rect 204382 313538 204466 313774
rect 204702 313538 240146 313774
rect 240382 313538 240466 313774
rect 240702 313538 276146 313774
rect 276382 313538 276466 313774
rect 276702 313538 312146 313774
rect 312382 313538 312466 313774
rect 312702 313538 348146 313774
rect 348382 313538 348466 313774
rect 348702 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 592650 313774
rect -8726 313454 592650 313538
rect -8726 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 24146 313454
rect 24382 313218 24466 313454
rect 24702 313218 60146 313454
rect 60382 313218 60466 313454
rect 60702 313218 96146 313454
rect 96382 313218 96466 313454
rect 96702 313218 132146 313454
rect 132382 313218 132466 313454
rect 132702 313218 168146 313454
rect 168382 313218 168466 313454
rect 168702 313218 204146 313454
rect 204382 313218 204466 313454
rect 204702 313218 240146 313454
rect 240382 313218 240466 313454
rect 240702 313218 276146 313454
rect 276382 313218 276466 313454
rect 276702 313218 312146 313454
rect 312382 313218 312466 313454
rect 312702 313218 348146 313454
rect 348382 313218 348466 313454
rect 348702 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 592650 313454
rect -8726 313186 592650 313218
rect -8726 310054 592650 310086
rect -8726 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 56426 310054
rect 56662 309818 56746 310054
rect 56982 309818 92426 310054
rect 92662 309818 92746 310054
rect 92982 309818 128426 310054
rect 128662 309818 128746 310054
rect 128982 309818 164426 310054
rect 164662 309818 164746 310054
rect 164982 309818 200426 310054
rect 200662 309818 200746 310054
rect 200982 309818 236426 310054
rect 236662 309818 236746 310054
rect 236982 309818 272426 310054
rect 272662 309818 272746 310054
rect 272982 309818 308426 310054
rect 308662 309818 308746 310054
rect 308982 309818 344426 310054
rect 344662 309818 344746 310054
rect 344982 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 592650 310054
rect -8726 309734 592650 309818
rect -8726 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 56426 309734
rect 56662 309498 56746 309734
rect 56982 309498 92426 309734
rect 92662 309498 92746 309734
rect 92982 309498 128426 309734
rect 128662 309498 128746 309734
rect 128982 309498 164426 309734
rect 164662 309498 164746 309734
rect 164982 309498 200426 309734
rect 200662 309498 200746 309734
rect 200982 309498 236426 309734
rect 236662 309498 236746 309734
rect 236982 309498 272426 309734
rect 272662 309498 272746 309734
rect 272982 309498 308426 309734
rect 308662 309498 308746 309734
rect 308982 309498 344426 309734
rect 344662 309498 344746 309734
rect 344982 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 592650 309734
rect -8726 309466 592650 309498
rect -8726 306334 592650 306366
rect -8726 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 52706 306334
rect 52942 306098 53026 306334
rect 53262 306098 88706 306334
rect 88942 306098 89026 306334
rect 89262 306098 124706 306334
rect 124942 306098 125026 306334
rect 125262 306098 160706 306334
rect 160942 306098 161026 306334
rect 161262 306098 196706 306334
rect 196942 306098 197026 306334
rect 197262 306098 232706 306334
rect 232942 306098 233026 306334
rect 233262 306098 268706 306334
rect 268942 306098 269026 306334
rect 269262 306098 304706 306334
rect 304942 306098 305026 306334
rect 305262 306098 340706 306334
rect 340942 306098 341026 306334
rect 341262 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 592650 306334
rect -8726 306014 592650 306098
rect -8726 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 52706 306014
rect 52942 305778 53026 306014
rect 53262 305778 88706 306014
rect 88942 305778 89026 306014
rect 89262 305778 124706 306014
rect 124942 305778 125026 306014
rect 125262 305778 160706 306014
rect 160942 305778 161026 306014
rect 161262 305778 196706 306014
rect 196942 305778 197026 306014
rect 197262 305778 232706 306014
rect 232942 305778 233026 306014
rect 233262 305778 268706 306014
rect 268942 305778 269026 306014
rect 269262 305778 304706 306014
rect 304942 305778 305026 306014
rect 305262 305778 340706 306014
rect 340942 305778 341026 306014
rect 341262 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 592650 306014
rect -8726 305746 592650 305778
rect -8726 302614 592650 302646
rect -8726 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 592650 302294
rect -8726 302026 592650 302058
rect -8726 298894 592650 298926
rect -8726 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 592650 298894
rect -8726 298574 592650 298658
rect -8726 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 592650 298574
rect -8726 298306 592650 298338
rect -8726 295174 592650 295206
rect -8726 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 592650 295174
rect -8726 294854 592650 294938
rect -8726 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 592650 294854
rect -8726 294586 592650 294618
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 281494 592650 281526
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 63866 281494
rect 64102 281258 64186 281494
rect 64422 281258 99866 281494
rect 100102 281258 100186 281494
rect 100422 281258 135866 281494
rect 136102 281258 136186 281494
rect 136422 281258 171866 281494
rect 172102 281258 172186 281494
rect 172422 281258 207866 281494
rect 208102 281258 208186 281494
rect 208422 281258 243866 281494
rect 244102 281258 244186 281494
rect 244422 281258 279866 281494
rect 280102 281258 280186 281494
rect 280422 281258 315866 281494
rect 316102 281258 316186 281494
rect 316422 281258 351866 281494
rect 352102 281258 352186 281494
rect 352422 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect -8726 281174 592650 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 63866 281174
rect 64102 280938 64186 281174
rect 64422 280938 99866 281174
rect 100102 280938 100186 281174
rect 100422 280938 135866 281174
rect 136102 280938 136186 281174
rect 136422 280938 171866 281174
rect 172102 280938 172186 281174
rect 172422 280938 207866 281174
rect 208102 280938 208186 281174
rect 208422 280938 243866 281174
rect 244102 280938 244186 281174
rect 244422 280938 279866 281174
rect 280102 280938 280186 281174
rect 280422 280938 315866 281174
rect 316102 280938 316186 281174
rect 316422 280938 351866 281174
rect 352102 280938 352186 281174
rect 352422 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect -8726 280906 592650 280938
rect -8726 277774 592650 277806
rect -8726 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 24146 277774
rect 24382 277538 24466 277774
rect 24702 277538 60146 277774
rect 60382 277538 60466 277774
rect 60702 277538 96146 277774
rect 96382 277538 96466 277774
rect 96702 277538 132146 277774
rect 132382 277538 132466 277774
rect 132702 277538 168146 277774
rect 168382 277538 168466 277774
rect 168702 277538 204146 277774
rect 204382 277538 204466 277774
rect 204702 277538 240146 277774
rect 240382 277538 240466 277774
rect 240702 277538 276146 277774
rect 276382 277538 276466 277774
rect 276702 277538 312146 277774
rect 312382 277538 312466 277774
rect 312702 277538 348146 277774
rect 348382 277538 348466 277774
rect 348702 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 592650 277774
rect -8726 277454 592650 277538
rect -8726 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 24146 277454
rect 24382 277218 24466 277454
rect 24702 277218 60146 277454
rect 60382 277218 60466 277454
rect 60702 277218 96146 277454
rect 96382 277218 96466 277454
rect 96702 277218 132146 277454
rect 132382 277218 132466 277454
rect 132702 277218 168146 277454
rect 168382 277218 168466 277454
rect 168702 277218 204146 277454
rect 204382 277218 204466 277454
rect 204702 277218 240146 277454
rect 240382 277218 240466 277454
rect 240702 277218 276146 277454
rect 276382 277218 276466 277454
rect 276702 277218 312146 277454
rect 312382 277218 312466 277454
rect 312702 277218 348146 277454
rect 348382 277218 348466 277454
rect 348702 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 592650 277454
rect -8726 277186 592650 277218
rect -8726 274054 592650 274086
rect -8726 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 56426 274054
rect 56662 273818 56746 274054
rect 56982 273818 92426 274054
rect 92662 273818 92746 274054
rect 92982 273818 128426 274054
rect 128662 273818 128746 274054
rect 128982 273818 164426 274054
rect 164662 273818 164746 274054
rect 164982 273818 200426 274054
rect 200662 273818 200746 274054
rect 200982 273818 236426 274054
rect 236662 273818 236746 274054
rect 236982 273818 272426 274054
rect 272662 273818 272746 274054
rect 272982 273818 308426 274054
rect 308662 273818 308746 274054
rect 308982 273818 344426 274054
rect 344662 273818 344746 274054
rect 344982 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 592650 274054
rect -8726 273734 592650 273818
rect -8726 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 56426 273734
rect 56662 273498 56746 273734
rect 56982 273498 92426 273734
rect 92662 273498 92746 273734
rect 92982 273498 128426 273734
rect 128662 273498 128746 273734
rect 128982 273498 164426 273734
rect 164662 273498 164746 273734
rect 164982 273498 200426 273734
rect 200662 273498 200746 273734
rect 200982 273498 236426 273734
rect 236662 273498 236746 273734
rect 236982 273498 272426 273734
rect 272662 273498 272746 273734
rect 272982 273498 308426 273734
rect 308662 273498 308746 273734
rect 308982 273498 344426 273734
rect 344662 273498 344746 273734
rect 344982 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 592650 273734
rect -8726 273466 592650 273498
rect -8726 270334 592650 270366
rect -8726 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 52706 270334
rect 52942 270098 53026 270334
rect 53262 270098 88706 270334
rect 88942 270098 89026 270334
rect 89262 270098 124706 270334
rect 124942 270098 125026 270334
rect 125262 270098 160706 270334
rect 160942 270098 161026 270334
rect 161262 270098 196706 270334
rect 196942 270098 197026 270334
rect 197262 270098 232706 270334
rect 232942 270098 233026 270334
rect 233262 270098 268706 270334
rect 268942 270098 269026 270334
rect 269262 270098 304706 270334
rect 304942 270098 305026 270334
rect 305262 270098 340706 270334
rect 340942 270098 341026 270334
rect 341262 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 592650 270334
rect -8726 270014 592650 270098
rect -8726 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 52706 270014
rect 52942 269778 53026 270014
rect 53262 269778 88706 270014
rect 88942 269778 89026 270014
rect 89262 269778 124706 270014
rect 124942 269778 125026 270014
rect 125262 269778 160706 270014
rect 160942 269778 161026 270014
rect 161262 269778 196706 270014
rect 196942 269778 197026 270014
rect 197262 269778 232706 270014
rect 232942 269778 233026 270014
rect 233262 269778 268706 270014
rect 268942 269778 269026 270014
rect 269262 269778 304706 270014
rect 304942 269778 305026 270014
rect 305262 269778 340706 270014
rect 340942 269778 341026 270014
rect 341262 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 592650 270014
rect -8726 269746 592650 269778
rect -8726 266614 592650 266646
rect -8726 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 592650 266294
rect -8726 266026 592650 266058
rect -8726 262894 592650 262926
rect -8726 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 592650 262894
rect -8726 262574 592650 262658
rect -8726 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 592650 262574
rect -8726 262306 592650 262338
rect -8726 259174 592650 259206
rect -8726 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 592650 259174
rect -8726 258854 592650 258938
rect -8726 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 592650 258854
rect -8726 258586 592650 258618
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 245494 592650 245526
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 63866 245494
rect 64102 245258 64186 245494
rect 64422 245258 99866 245494
rect 100102 245258 100186 245494
rect 100422 245258 135866 245494
rect 136102 245258 136186 245494
rect 136422 245258 171866 245494
rect 172102 245258 172186 245494
rect 172422 245258 207866 245494
rect 208102 245258 208186 245494
rect 208422 245258 243866 245494
rect 244102 245258 244186 245494
rect 244422 245258 279866 245494
rect 280102 245258 280186 245494
rect 280422 245258 315866 245494
rect 316102 245258 316186 245494
rect 316422 245258 351866 245494
rect 352102 245258 352186 245494
rect 352422 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 495866 245494
rect 496102 245258 496186 245494
rect 496422 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect -8726 245174 592650 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 63866 245174
rect 64102 244938 64186 245174
rect 64422 244938 99866 245174
rect 100102 244938 100186 245174
rect 100422 244938 135866 245174
rect 136102 244938 136186 245174
rect 136422 244938 171866 245174
rect 172102 244938 172186 245174
rect 172422 244938 207866 245174
rect 208102 244938 208186 245174
rect 208422 244938 243866 245174
rect 244102 244938 244186 245174
rect 244422 244938 279866 245174
rect 280102 244938 280186 245174
rect 280422 244938 315866 245174
rect 316102 244938 316186 245174
rect 316422 244938 351866 245174
rect 352102 244938 352186 245174
rect 352422 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 495866 245174
rect 496102 244938 496186 245174
rect 496422 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect -8726 244906 592650 244938
rect -8726 241774 592650 241806
rect -8726 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 24146 241774
rect 24382 241538 24466 241774
rect 24702 241538 60146 241774
rect 60382 241538 60466 241774
rect 60702 241538 96146 241774
rect 96382 241538 96466 241774
rect 96702 241538 132146 241774
rect 132382 241538 132466 241774
rect 132702 241538 168146 241774
rect 168382 241538 168466 241774
rect 168702 241538 204146 241774
rect 204382 241538 204466 241774
rect 204702 241538 240146 241774
rect 240382 241538 240466 241774
rect 240702 241538 276146 241774
rect 276382 241538 276466 241774
rect 276702 241538 312146 241774
rect 312382 241538 312466 241774
rect 312702 241538 348146 241774
rect 348382 241538 348466 241774
rect 348702 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 492146 241774
rect 492382 241538 492466 241774
rect 492702 241538 528146 241774
rect 528382 241538 528466 241774
rect 528702 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 592650 241774
rect -8726 241454 592650 241538
rect -8726 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 24146 241454
rect 24382 241218 24466 241454
rect 24702 241218 60146 241454
rect 60382 241218 60466 241454
rect 60702 241218 96146 241454
rect 96382 241218 96466 241454
rect 96702 241218 132146 241454
rect 132382 241218 132466 241454
rect 132702 241218 168146 241454
rect 168382 241218 168466 241454
rect 168702 241218 204146 241454
rect 204382 241218 204466 241454
rect 204702 241218 240146 241454
rect 240382 241218 240466 241454
rect 240702 241218 276146 241454
rect 276382 241218 276466 241454
rect 276702 241218 312146 241454
rect 312382 241218 312466 241454
rect 312702 241218 348146 241454
rect 348382 241218 348466 241454
rect 348702 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 492146 241454
rect 492382 241218 492466 241454
rect 492702 241218 528146 241454
rect 528382 241218 528466 241454
rect 528702 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 592650 241454
rect -8726 241186 592650 241218
rect -8726 238054 592650 238086
rect -8726 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 56426 238054
rect 56662 237818 56746 238054
rect 56982 237818 128426 238054
rect 128662 237818 128746 238054
rect 128982 237818 164426 238054
rect 164662 237818 164746 238054
rect 164982 237818 200426 238054
rect 200662 237818 200746 238054
rect 200982 237818 236426 238054
rect 236662 237818 236746 238054
rect 236982 237818 272426 238054
rect 272662 237818 272746 238054
rect 272982 237818 308426 238054
rect 308662 237818 308746 238054
rect 308982 237818 344426 238054
rect 344662 237818 344746 238054
rect 344982 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 488426 238054
rect 488662 237818 488746 238054
rect 488982 237818 524426 238054
rect 524662 237818 524746 238054
rect 524982 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 592650 238054
rect -8726 237734 592650 237818
rect -8726 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 56426 237734
rect 56662 237498 56746 237734
rect 56982 237498 128426 237734
rect 128662 237498 128746 237734
rect 128982 237498 164426 237734
rect 164662 237498 164746 237734
rect 164982 237498 200426 237734
rect 200662 237498 200746 237734
rect 200982 237498 236426 237734
rect 236662 237498 236746 237734
rect 236982 237498 272426 237734
rect 272662 237498 272746 237734
rect 272982 237498 308426 237734
rect 308662 237498 308746 237734
rect 308982 237498 344426 237734
rect 344662 237498 344746 237734
rect 344982 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 488426 237734
rect 488662 237498 488746 237734
rect 488982 237498 524426 237734
rect 524662 237498 524746 237734
rect 524982 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 592650 237734
rect -8726 237466 592650 237498
rect -8726 234334 592650 234366
rect -8726 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 52706 234334
rect 52942 234098 53026 234334
rect 53262 234098 124706 234334
rect 124942 234098 125026 234334
rect 125262 234098 160706 234334
rect 160942 234098 161026 234334
rect 161262 234098 196706 234334
rect 196942 234098 197026 234334
rect 197262 234098 232706 234334
rect 232942 234098 233026 234334
rect 233262 234098 268706 234334
rect 268942 234098 269026 234334
rect 269262 234098 304706 234334
rect 304942 234098 305026 234334
rect 305262 234098 340706 234334
rect 340942 234098 341026 234334
rect 341262 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 484706 234334
rect 484942 234098 485026 234334
rect 485262 234098 520706 234334
rect 520942 234098 521026 234334
rect 521262 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 592650 234334
rect -8726 234014 592650 234098
rect -8726 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 52706 234014
rect 52942 233778 53026 234014
rect 53262 233778 124706 234014
rect 124942 233778 125026 234014
rect 125262 233778 160706 234014
rect 160942 233778 161026 234014
rect 161262 233778 196706 234014
rect 196942 233778 197026 234014
rect 197262 233778 232706 234014
rect 232942 233778 233026 234014
rect 233262 233778 268706 234014
rect 268942 233778 269026 234014
rect 269262 233778 304706 234014
rect 304942 233778 305026 234014
rect 305262 233778 340706 234014
rect 340942 233778 341026 234014
rect 341262 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 484706 234014
rect 484942 233778 485026 234014
rect 485262 233778 520706 234014
rect 520942 233778 521026 234014
rect 521262 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 592650 234014
rect -8726 233746 592650 233778
rect -8726 230614 592650 230646
rect -8726 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 592650 230294
rect -8726 230026 592650 230058
rect -8726 226894 592650 226926
rect -8726 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 592650 226894
rect -8726 226574 592650 226658
rect -8726 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 592650 226574
rect -8726 226306 592650 226338
rect -8726 223174 592650 223206
rect -8726 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 89610 223174
rect 89846 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 189610 223174
rect 189846 222938 220330 223174
rect 220566 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 592650 223174
rect -8726 222854 592650 222938
rect -8726 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 89610 222854
rect 89846 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 189610 222854
rect 189846 222618 220330 222854
rect 220566 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 592650 222854
rect -8726 222586 592650 222618
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 74250 219454
rect 74486 219218 104970 219454
rect 105206 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 174250 219454
rect 174486 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 204970 219454
rect 205206 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 74250 219134
rect 74486 218898 104970 219134
rect 105206 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 174250 219134
rect 174486 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 204970 219134
rect 205206 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 209494 592650 209526
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 63866 209494
rect 64102 209258 64186 209494
rect 64422 209258 99866 209494
rect 100102 209258 100186 209494
rect 100422 209258 135866 209494
rect 136102 209258 136186 209494
rect 136422 209258 171866 209494
rect 172102 209258 172186 209494
rect 172422 209258 243866 209494
rect 244102 209258 244186 209494
rect 244422 209258 279866 209494
rect 280102 209258 280186 209494
rect 280422 209258 315866 209494
rect 316102 209258 316186 209494
rect 316422 209258 351866 209494
rect 352102 209258 352186 209494
rect 352422 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 495866 209494
rect 496102 209258 496186 209494
rect 496422 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect -8726 209174 592650 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 63866 209174
rect 64102 208938 64186 209174
rect 64422 208938 99866 209174
rect 100102 208938 100186 209174
rect 100422 208938 135866 209174
rect 136102 208938 136186 209174
rect 136422 208938 171866 209174
rect 172102 208938 172186 209174
rect 172422 208938 243866 209174
rect 244102 208938 244186 209174
rect 244422 208938 279866 209174
rect 280102 208938 280186 209174
rect 280422 208938 315866 209174
rect 316102 208938 316186 209174
rect 316422 208938 351866 209174
rect 352102 208938 352186 209174
rect 352422 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 495866 209174
rect 496102 208938 496186 209174
rect 496422 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect -8726 208906 592650 208938
rect -8726 205774 592650 205806
rect -8726 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 24146 205774
rect 24382 205538 24466 205774
rect 24702 205538 60146 205774
rect 60382 205538 60466 205774
rect 60702 205538 96146 205774
rect 96382 205538 96466 205774
rect 96702 205538 132146 205774
rect 132382 205538 132466 205774
rect 132702 205538 168146 205774
rect 168382 205538 168466 205774
rect 168702 205538 240146 205774
rect 240382 205538 240466 205774
rect 240702 205538 276146 205774
rect 276382 205538 276466 205774
rect 276702 205538 312146 205774
rect 312382 205538 312466 205774
rect 312702 205538 348146 205774
rect 348382 205538 348466 205774
rect 348702 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 420146 205774
rect 420382 205538 420466 205774
rect 420702 205538 456146 205774
rect 456382 205538 456466 205774
rect 456702 205538 492146 205774
rect 492382 205538 492466 205774
rect 492702 205538 528146 205774
rect 528382 205538 528466 205774
rect 528702 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 592650 205774
rect -8726 205454 592650 205538
rect -8726 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 24146 205454
rect 24382 205218 24466 205454
rect 24702 205218 60146 205454
rect 60382 205218 60466 205454
rect 60702 205218 96146 205454
rect 96382 205218 96466 205454
rect 96702 205218 132146 205454
rect 132382 205218 132466 205454
rect 132702 205218 168146 205454
rect 168382 205218 168466 205454
rect 168702 205218 240146 205454
rect 240382 205218 240466 205454
rect 240702 205218 276146 205454
rect 276382 205218 276466 205454
rect 276702 205218 312146 205454
rect 312382 205218 312466 205454
rect 312702 205218 348146 205454
rect 348382 205218 348466 205454
rect 348702 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 420146 205454
rect 420382 205218 420466 205454
rect 420702 205218 456146 205454
rect 456382 205218 456466 205454
rect 456702 205218 492146 205454
rect 492382 205218 492466 205454
rect 492702 205218 528146 205454
rect 528382 205218 528466 205454
rect 528702 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 592650 205454
rect -8726 205186 592650 205218
rect -8726 202054 592650 202086
rect -8726 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 56426 202054
rect 56662 201818 56746 202054
rect 56982 201818 92426 202054
rect 92662 201818 92746 202054
rect 92982 201818 128426 202054
rect 128662 201818 128746 202054
rect 128982 201818 164426 202054
rect 164662 201818 164746 202054
rect 164982 201818 236426 202054
rect 236662 201818 236746 202054
rect 236982 201818 272426 202054
rect 272662 201818 272746 202054
rect 272982 201818 308426 202054
rect 308662 201818 308746 202054
rect 308982 201818 344426 202054
rect 344662 201818 344746 202054
rect 344982 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 488426 202054
rect 488662 201818 488746 202054
rect 488982 201818 524426 202054
rect 524662 201818 524746 202054
rect 524982 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 592650 202054
rect -8726 201734 592650 201818
rect -8726 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 56426 201734
rect 56662 201498 56746 201734
rect 56982 201498 92426 201734
rect 92662 201498 92746 201734
rect 92982 201498 128426 201734
rect 128662 201498 128746 201734
rect 128982 201498 164426 201734
rect 164662 201498 164746 201734
rect 164982 201498 236426 201734
rect 236662 201498 236746 201734
rect 236982 201498 272426 201734
rect 272662 201498 272746 201734
rect 272982 201498 308426 201734
rect 308662 201498 308746 201734
rect 308982 201498 344426 201734
rect 344662 201498 344746 201734
rect 344982 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 488426 201734
rect 488662 201498 488746 201734
rect 488982 201498 524426 201734
rect 524662 201498 524746 201734
rect 524982 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 592650 201734
rect -8726 201466 592650 201498
rect -8726 198334 592650 198366
rect -8726 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 52706 198334
rect 52942 198098 53026 198334
rect 53262 198098 88706 198334
rect 88942 198098 89026 198334
rect 89262 198098 124706 198334
rect 124942 198098 125026 198334
rect 125262 198098 160706 198334
rect 160942 198098 161026 198334
rect 161262 198098 232706 198334
rect 232942 198098 233026 198334
rect 233262 198098 268706 198334
rect 268942 198098 269026 198334
rect 269262 198098 304706 198334
rect 304942 198098 305026 198334
rect 305262 198098 340706 198334
rect 340942 198098 341026 198334
rect 341262 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 592650 198334
rect -8726 198014 592650 198098
rect -8726 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 52706 198014
rect 52942 197778 53026 198014
rect 53262 197778 88706 198014
rect 88942 197778 89026 198014
rect 89262 197778 124706 198014
rect 124942 197778 125026 198014
rect 125262 197778 160706 198014
rect 160942 197778 161026 198014
rect 161262 197778 232706 198014
rect 232942 197778 233026 198014
rect 233262 197778 268706 198014
rect 268942 197778 269026 198014
rect 269262 197778 304706 198014
rect 304942 197778 305026 198014
rect 305262 197778 340706 198014
rect 340942 197778 341026 198014
rect 341262 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 592650 198014
rect -8726 197746 592650 197778
rect -8726 194614 592650 194646
rect -8726 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 592650 194294
rect -8726 194026 592650 194058
rect -8726 190894 592650 190926
rect -8726 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 592650 190894
rect -8726 190574 592650 190658
rect -8726 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 592650 190574
rect -8726 190306 592650 190338
rect -8726 187174 592650 187206
rect -8726 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 189610 187174
rect 189846 186938 220330 187174
rect 220566 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 592650 187174
rect -8726 186854 592650 186938
rect -8726 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 189610 186854
rect 189846 186618 220330 186854
rect 220566 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 592650 186854
rect -8726 186586 592650 186618
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 174250 183454
rect 174486 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 204970 183454
rect 205206 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 174250 183134
rect 174486 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 204970 183134
rect 205206 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 173494 592650 173526
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 63866 173494
rect 64102 173258 64186 173494
rect 64422 173258 99866 173494
rect 100102 173258 100186 173494
rect 100422 173258 135866 173494
rect 136102 173258 136186 173494
rect 136422 173258 171866 173494
rect 172102 173258 172186 173494
rect 172422 173258 207866 173494
rect 208102 173258 208186 173494
rect 208422 173258 243866 173494
rect 244102 173258 244186 173494
rect 244422 173258 279866 173494
rect 280102 173258 280186 173494
rect 280422 173258 315866 173494
rect 316102 173258 316186 173494
rect 316422 173258 351866 173494
rect 352102 173258 352186 173494
rect 352422 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 495866 173494
rect 496102 173258 496186 173494
rect 496422 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect -8726 173174 592650 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 63866 173174
rect 64102 172938 64186 173174
rect 64422 172938 99866 173174
rect 100102 172938 100186 173174
rect 100422 172938 135866 173174
rect 136102 172938 136186 173174
rect 136422 172938 171866 173174
rect 172102 172938 172186 173174
rect 172422 172938 207866 173174
rect 208102 172938 208186 173174
rect 208422 172938 243866 173174
rect 244102 172938 244186 173174
rect 244422 172938 279866 173174
rect 280102 172938 280186 173174
rect 280422 172938 315866 173174
rect 316102 172938 316186 173174
rect 316422 172938 351866 173174
rect 352102 172938 352186 173174
rect 352422 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 495866 173174
rect 496102 172938 496186 173174
rect 496422 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect -8726 172906 592650 172938
rect -8726 169774 592650 169806
rect -8726 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 24146 169774
rect 24382 169538 24466 169774
rect 24702 169538 60146 169774
rect 60382 169538 60466 169774
rect 60702 169538 96146 169774
rect 96382 169538 96466 169774
rect 96702 169538 132146 169774
rect 132382 169538 132466 169774
rect 132702 169538 168146 169774
rect 168382 169538 168466 169774
rect 168702 169538 204146 169774
rect 204382 169538 204466 169774
rect 204702 169538 240146 169774
rect 240382 169538 240466 169774
rect 240702 169538 276146 169774
rect 276382 169538 276466 169774
rect 276702 169538 312146 169774
rect 312382 169538 312466 169774
rect 312702 169538 348146 169774
rect 348382 169538 348466 169774
rect 348702 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 420146 169774
rect 420382 169538 420466 169774
rect 420702 169538 456146 169774
rect 456382 169538 456466 169774
rect 456702 169538 492146 169774
rect 492382 169538 492466 169774
rect 492702 169538 528146 169774
rect 528382 169538 528466 169774
rect 528702 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 592650 169774
rect -8726 169454 592650 169538
rect -8726 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 24146 169454
rect 24382 169218 24466 169454
rect 24702 169218 60146 169454
rect 60382 169218 60466 169454
rect 60702 169218 96146 169454
rect 96382 169218 96466 169454
rect 96702 169218 132146 169454
rect 132382 169218 132466 169454
rect 132702 169218 168146 169454
rect 168382 169218 168466 169454
rect 168702 169218 204146 169454
rect 204382 169218 204466 169454
rect 204702 169218 240146 169454
rect 240382 169218 240466 169454
rect 240702 169218 276146 169454
rect 276382 169218 276466 169454
rect 276702 169218 312146 169454
rect 312382 169218 312466 169454
rect 312702 169218 348146 169454
rect 348382 169218 348466 169454
rect 348702 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 420146 169454
rect 420382 169218 420466 169454
rect 420702 169218 456146 169454
rect 456382 169218 456466 169454
rect 456702 169218 492146 169454
rect 492382 169218 492466 169454
rect 492702 169218 528146 169454
rect 528382 169218 528466 169454
rect 528702 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 592650 169454
rect -8726 169186 592650 169218
rect -8726 166054 592650 166086
rect -8726 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 56426 166054
rect 56662 165818 56746 166054
rect 56982 165818 92426 166054
rect 92662 165818 92746 166054
rect 92982 165818 128426 166054
rect 128662 165818 128746 166054
rect 128982 165818 164426 166054
rect 164662 165818 164746 166054
rect 164982 165818 200426 166054
rect 200662 165818 200746 166054
rect 200982 165818 236426 166054
rect 236662 165818 236746 166054
rect 236982 165818 272426 166054
rect 272662 165818 272746 166054
rect 272982 165818 308426 166054
rect 308662 165818 308746 166054
rect 308982 165818 344426 166054
rect 344662 165818 344746 166054
rect 344982 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 592650 166054
rect -8726 165734 592650 165818
rect -8726 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 56426 165734
rect 56662 165498 56746 165734
rect 56982 165498 92426 165734
rect 92662 165498 92746 165734
rect 92982 165498 128426 165734
rect 128662 165498 128746 165734
rect 128982 165498 164426 165734
rect 164662 165498 164746 165734
rect 164982 165498 200426 165734
rect 200662 165498 200746 165734
rect 200982 165498 236426 165734
rect 236662 165498 236746 165734
rect 236982 165498 272426 165734
rect 272662 165498 272746 165734
rect 272982 165498 308426 165734
rect 308662 165498 308746 165734
rect 308982 165498 344426 165734
rect 344662 165498 344746 165734
rect 344982 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 592650 165734
rect -8726 165466 592650 165498
rect -8726 162334 592650 162366
rect -8726 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 52706 162334
rect 52942 162098 53026 162334
rect 53262 162098 88706 162334
rect 88942 162098 89026 162334
rect 89262 162098 124706 162334
rect 124942 162098 125026 162334
rect 125262 162098 160706 162334
rect 160942 162098 161026 162334
rect 161262 162098 196706 162334
rect 196942 162098 197026 162334
rect 197262 162098 232706 162334
rect 232942 162098 233026 162334
rect 233262 162098 268706 162334
rect 268942 162098 269026 162334
rect 269262 162098 304706 162334
rect 304942 162098 305026 162334
rect 305262 162098 340706 162334
rect 340942 162098 341026 162334
rect 341262 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 448706 162334
rect 448942 162098 449026 162334
rect 449262 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 592650 162334
rect -8726 162014 592650 162098
rect -8726 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 52706 162014
rect 52942 161778 53026 162014
rect 53262 161778 88706 162014
rect 88942 161778 89026 162014
rect 89262 161778 124706 162014
rect 124942 161778 125026 162014
rect 125262 161778 160706 162014
rect 160942 161778 161026 162014
rect 161262 161778 196706 162014
rect 196942 161778 197026 162014
rect 197262 161778 232706 162014
rect 232942 161778 233026 162014
rect 233262 161778 268706 162014
rect 268942 161778 269026 162014
rect 269262 161778 304706 162014
rect 304942 161778 305026 162014
rect 305262 161778 340706 162014
rect 340942 161778 341026 162014
rect 341262 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 448706 162014
rect 448942 161778 449026 162014
rect 449262 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 592650 162014
rect -8726 161746 592650 161778
rect -8726 158614 592650 158646
rect -8726 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 592650 158294
rect -8726 158026 592650 158058
rect -8726 154894 592650 154926
rect -8726 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 592650 154894
rect -8726 154574 592650 154658
rect -8726 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 592650 154574
rect -8726 154306 592650 154338
rect -8726 151174 592650 151206
rect -8726 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 592650 151174
rect -8726 150854 592650 150938
rect -8726 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 592650 150854
rect -8726 150586 592650 150618
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 137494 592650 137526
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 63866 137494
rect 64102 137258 64186 137494
rect 64422 137258 99866 137494
rect 100102 137258 100186 137494
rect 100422 137258 135866 137494
rect 136102 137258 136186 137494
rect 136422 137258 171866 137494
rect 172102 137258 172186 137494
rect 172422 137258 207866 137494
rect 208102 137258 208186 137494
rect 208422 137258 243866 137494
rect 244102 137258 244186 137494
rect 244422 137258 279866 137494
rect 280102 137258 280186 137494
rect 280422 137258 315866 137494
rect 316102 137258 316186 137494
rect 316422 137258 351866 137494
rect 352102 137258 352186 137494
rect 352422 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 423866 137494
rect 424102 137258 424186 137494
rect 424422 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 495866 137494
rect 496102 137258 496186 137494
rect 496422 137258 531866 137494
rect 532102 137258 532186 137494
rect 532422 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect -8726 137174 592650 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 63866 137174
rect 64102 136938 64186 137174
rect 64422 136938 99866 137174
rect 100102 136938 100186 137174
rect 100422 136938 135866 137174
rect 136102 136938 136186 137174
rect 136422 136938 171866 137174
rect 172102 136938 172186 137174
rect 172422 136938 207866 137174
rect 208102 136938 208186 137174
rect 208422 136938 243866 137174
rect 244102 136938 244186 137174
rect 244422 136938 279866 137174
rect 280102 136938 280186 137174
rect 280422 136938 315866 137174
rect 316102 136938 316186 137174
rect 316422 136938 351866 137174
rect 352102 136938 352186 137174
rect 352422 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 423866 137174
rect 424102 136938 424186 137174
rect 424422 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 495866 137174
rect 496102 136938 496186 137174
rect 496422 136938 531866 137174
rect 532102 136938 532186 137174
rect 532422 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect -8726 136906 592650 136938
rect -8726 133774 592650 133806
rect -8726 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 24146 133774
rect 24382 133538 24466 133774
rect 24702 133538 60146 133774
rect 60382 133538 60466 133774
rect 60702 133538 96146 133774
rect 96382 133538 96466 133774
rect 96702 133538 132146 133774
rect 132382 133538 132466 133774
rect 132702 133538 168146 133774
rect 168382 133538 168466 133774
rect 168702 133538 204146 133774
rect 204382 133538 204466 133774
rect 204702 133538 240146 133774
rect 240382 133538 240466 133774
rect 240702 133538 276146 133774
rect 276382 133538 276466 133774
rect 276702 133538 312146 133774
rect 312382 133538 312466 133774
rect 312702 133538 348146 133774
rect 348382 133538 348466 133774
rect 348702 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 420146 133774
rect 420382 133538 420466 133774
rect 420702 133538 456146 133774
rect 456382 133538 456466 133774
rect 456702 133538 492146 133774
rect 492382 133538 492466 133774
rect 492702 133538 528146 133774
rect 528382 133538 528466 133774
rect 528702 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 592650 133774
rect -8726 133454 592650 133538
rect -8726 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 24146 133454
rect 24382 133218 24466 133454
rect 24702 133218 60146 133454
rect 60382 133218 60466 133454
rect 60702 133218 96146 133454
rect 96382 133218 96466 133454
rect 96702 133218 132146 133454
rect 132382 133218 132466 133454
rect 132702 133218 168146 133454
rect 168382 133218 168466 133454
rect 168702 133218 204146 133454
rect 204382 133218 204466 133454
rect 204702 133218 240146 133454
rect 240382 133218 240466 133454
rect 240702 133218 276146 133454
rect 276382 133218 276466 133454
rect 276702 133218 312146 133454
rect 312382 133218 312466 133454
rect 312702 133218 348146 133454
rect 348382 133218 348466 133454
rect 348702 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 420146 133454
rect 420382 133218 420466 133454
rect 420702 133218 456146 133454
rect 456382 133218 456466 133454
rect 456702 133218 492146 133454
rect 492382 133218 492466 133454
rect 492702 133218 528146 133454
rect 528382 133218 528466 133454
rect 528702 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 592650 133454
rect -8726 133186 592650 133218
rect -8726 130054 592650 130086
rect -8726 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 56426 130054
rect 56662 129818 56746 130054
rect 56982 129818 92426 130054
rect 92662 129818 92746 130054
rect 92982 129818 128426 130054
rect 128662 129818 128746 130054
rect 128982 129818 164426 130054
rect 164662 129818 164746 130054
rect 164982 129818 200426 130054
rect 200662 129818 200746 130054
rect 200982 129818 236426 130054
rect 236662 129818 236746 130054
rect 236982 129818 272426 130054
rect 272662 129818 272746 130054
rect 272982 129818 308426 130054
rect 308662 129818 308746 130054
rect 308982 129818 344426 130054
rect 344662 129818 344746 130054
rect 344982 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 416426 130054
rect 416662 129818 416746 130054
rect 416982 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 488426 130054
rect 488662 129818 488746 130054
rect 488982 129818 524426 130054
rect 524662 129818 524746 130054
rect 524982 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 592650 130054
rect -8726 129734 592650 129818
rect -8726 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 56426 129734
rect 56662 129498 56746 129734
rect 56982 129498 92426 129734
rect 92662 129498 92746 129734
rect 92982 129498 128426 129734
rect 128662 129498 128746 129734
rect 128982 129498 164426 129734
rect 164662 129498 164746 129734
rect 164982 129498 200426 129734
rect 200662 129498 200746 129734
rect 200982 129498 236426 129734
rect 236662 129498 236746 129734
rect 236982 129498 272426 129734
rect 272662 129498 272746 129734
rect 272982 129498 308426 129734
rect 308662 129498 308746 129734
rect 308982 129498 344426 129734
rect 344662 129498 344746 129734
rect 344982 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 416426 129734
rect 416662 129498 416746 129734
rect 416982 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 488426 129734
rect 488662 129498 488746 129734
rect 488982 129498 524426 129734
rect 524662 129498 524746 129734
rect 524982 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 592650 129734
rect -8726 129466 592650 129498
rect -8726 126334 592650 126366
rect -8726 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 52706 126334
rect 52942 126098 53026 126334
rect 53262 126098 88706 126334
rect 88942 126098 89026 126334
rect 89262 126098 124706 126334
rect 124942 126098 125026 126334
rect 125262 126098 160706 126334
rect 160942 126098 161026 126334
rect 161262 126098 196706 126334
rect 196942 126098 197026 126334
rect 197262 126098 232706 126334
rect 232942 126098 233026 126334
rect 233262 126098 268706 126334
rect 268942 126098 269026 126334
rect 269262 126098 304706 126334
rect 304942 126098 305026 126334
rect 305262 126098 340706 126334
rect 340942 126098 341026 126334
rect 341262 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 448706 126334
rect 448942 126098 449026 126334
rect 449262 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 520706 126334
rect 520942 126098 521026 126334
rect 521262 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 592650 126334
rect -8726 126014 592650 126098
rect -8726 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 52706 126014
rect 52942 125778 53026 126014
rect 53262 125778 88706 126014
rect 88942 125778 89026 126014
rect 89262 125778 124706 126014
rect 124942 125778 125026 126014
rect 125262 125778 160706 126014
rect 160942 125778 161026 126014
rect 161262 125778 196706 126014
rect 196942 125778 197026 126014
rect 197262 125778 232706 126014
rect 232942 125778 233026 126014
rect 233262 125778 268706 126014
rect 268942 125778 269026 126014
rect 269262 125778 304706 126014
rect 304942 125778 305026 126014
rect 305262 125778 340706 126014
rect 340942 125778 341026 126014
rect 341262 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 448706 126014
rect 448942 125778 449026 126014
rect 449262 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 520706 126014
rect 520942 125778 521026 126014
rect 521262 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 592650 126014
rect -8726 125746 592650 125778
rect -8726 122614 592650 122646
rect -8726 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 592650 122294
rect -8726 122026 592650 122058
rect -8726 118894 592650 118926
rect -8726 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 592650 118894
rect -8726 118574 592650 118658
rect -8726 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 592650 118574
rect -8726 118306 592650 118338
rect -8726 115174 592650 115206
rect -8726 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 177932 115174
rect 178168 114938 184878 115174
rect 185114 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 191824 115174
rect 192060 114938 198770 115174
rect 199006 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 592650 115174
rect -8726 114854 592650 114938
rect -8726 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 177932 114854
rect 178168 114618 184878 114854
rect 185114 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 191824 114854
rect 192060 114618 198770 114854
rect 199006 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 592650 114854
rect -8726 114586 592650 114618
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 174459 111454
rect 174695 111218 181405 111454
rect 181641 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 188351 111454
rect 188587 111218 195297 111454
rect 195533 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 174459 111134
rect 174695 110898 181405 111134
rect 181641 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 188351 111134
rect 188587 110898 195297 111134
rect 195533 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 101494 592650 101526
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 63866 101494
rect 64102 101258 64186 101494
rect 64422 101258 135866 101494
rect 136102 101258 136186 101494
rect 136422 101258 171866 101494
rect 172102 101258 172186 101494
rect 172422 101258 207866 101494
rect 208102 101258 208186 101494
rect 208422 101258 243866 101494
rect 244102 101258 244186 101494
rect 244422 101258 279866 101494
rect 280102 101258 280186 101494
rect 280422 101258 315866 101494
rect 316102 101258 316186 101494
rect 316422 101258 351866 101494
rect 352102 101258 352186 101494
rect 352422 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 495866 101494
rect 496102 101258 496186 101494
rect 496422 101258 531866 101494
rect 532102 101258 532186 101494
rect 532422 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect -8726 101174 592650 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 63866 101174
rect 64102 100938 64186 101174
rect 64422 100938 135866 101174
rect 136102 100938 136186 101174
rect 136422 100938 171866 101174
rect 172102 100938 172186 101174
rect 172422 100938 207866 101174
rect 208102 100938 208186 101174
rect 208422 100938 243866 101174
rect 244102 100938 244186 101174
rect 244422 100938 279866 101174
rect 280102 100938 280186 101174
rect 280422 100938 315866 101174
rect 316102 100938 316186 101174
rect 316422 100938 351866 101174
rect 352102 100938 352186 101174
rect 352422 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 495866 101174
rect 496102 100938 496186 101174
rect 496422 100938 531866 101174
rect 532102 100938 532186 101174
rect 532422 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect -8726 100906 592650 100938
rect -8726 97774 592650 97806
rect -8726 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 24146 97774
rect 24382 97538 24466 97774
rect 24702 97538 60146 97774
rect 60382 97538 60466 97774
rect 60702 97538 132146 97774
rect 132382 97538 132466 97774
rect 132702 97538 168146 97774
rect 168382 97538 168466 97774
rect 168702 97538 204146 97774
rect 204382 97538 204466 97774
rect 204702 97538 240146 97774
rect 240382 97538 240466 97774
rect 240702 97538 276146 97774
rect 276382 97538 276466 97774
rect 276702 97538 312146 97774
rect 312382 97538 312466 97774
rect 312702 97538 348146 97774
rect 348382 97538 348466 97774
rect 348702 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 420146 97774
rect 420382 97538 420466 97774
rect 420702 97538 456146 97774
rect 456382 97538 456466 97774
rect 456702 97538 492146 97774
rect 492382 97538 492466 97774
rect 492702 97538 528146 97774
rect 528382 97538 528466 97774
rect 528702 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 592650 97774
rect -8726 97454 592650 97538
rect -8726 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 24146 97454
rect 24382 97218 24466 97454
rect 24702 97218 60146 97454
rect 60382 97218 60466 97454
rect 60702 97218 132146 97454
rect 132382 97218 132466 97454
rect 132702 97218 168146 97454
rect 168382 97218 168466 97454
rect 168702 97218 204146 97454
rect 204382 97218 204466 97454
rect 204702 97218 240146 97454
rect 240382 97218 240466 97454
rect 240702 97218 276146 97454
rect 276382 97218 276466 97454
rect 276702 97218 312146 97454
rect 312382 97218 312466 97454
rect 312702 97218 348146 97454
rect 348382 97218 348466 97454
rect 348702 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 420146 97454
rect 420382 97218 420466 97454
rect 420702 97218 456146 97454
rect 456382 97218 456466 97454
rect 456702 97218 492146 97454
rect 492382 97218 492466 97454
rect 492702 97218 528146 97454
rect 528382 97218 528466 97454
rect 528702 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 592650 97454
rect -8726 97186 592650 97218
rect -8726 94054 592650 94086
rect -8726 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 56426 94054
rect 56662 93818 56746 94054
rect 56982 93818 128426 94054
rect 128662 93818 128746 94054
rect 128982 93818 164426 94054
rect 164662 93818 164746 94054
rect 164982 93818 200426 94054
rect 200662 93818 200746 94054
rect 200982 93818 236426 94054
rect 236662 93818 236746 94054
rect 236982 93818 272426 94054
rect 272662 93818 272746 94054
rect 272982 93818 308426 94054
rect 308662 93818 308746 94054
rect 308982 93818 344426 94054
rect 344662 93818 344746 94054
rect 344982 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 488426 94054
rect 488662 93818 488746 94054
rect 488982 93818 524426 94054
rect 524662 93818 524746 94054
rect 524982 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 592650 94054
rect -8726 93734 592650 93818
rect -8726 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 56426 93734
rect 56662 93498 56746 93734
rect 56982 93498 128426 93734
rect 128662 93498 128746 93734
rect 128982 93498 164426 93734
rect 164662 93498 164746 93734
rect 164982 93498 200426 93734
rect 200662 93498 200746 93734
rect 200982 93498 236426 93734
rect 236662 93498 236746 93734
rect 236982 93498 272426 93734
rect 272662 93498 272746 93734
rect 272982 93498 308426 93734
rect 308662 93498 308746 93734
rect 308982 93498 344426 93734
rect 344662 93498 344746 93734
rect 344982 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 488426 93734
rect 488662 93498 488746 93734
rect 488982 93498 524426 93734
rect 524662 93498 524746 93734
rect 524982 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 592650 93734
rect -8726 93466 592650 93498
rect -8726 90334 592650 90366
rect -8726 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 52706 90334
rect 52942 90098 53026 90334
rect 53262 90098 88706 90334
rect 88942 90098 89026 90334
rect 89262 90098 124706 90334
rect 124942 90098 125026 90334
rect 125262 90098 160706 90334
rect 160942 90098 161026 90334
rect 161262 90098 196706 90334
rect 196942 90098 197026 90334
rect 197262 90098 232706 90334
rect 232942 90098 233026 90334
rect 233262 90098 268706 90334
rect 268942 90098 269026 90334
rect 269262 90098 304706 90334
rect 304942 90098 305026 90334
rect 305262 90098 340706 90334
rect 340942 90098 341026 90334
rect 341262 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 412706 90334
rect 412942 90098 413026 90334
rect 413262 90098 448706 90334
rect 448942 90098 449026 90334
rect 449262 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 520706 90334
rect 520942 90098 521026 90334
rect 521262 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 592650 90334
rect -8726 90014 592650 90098
rect -8726 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 52706 90014
rect 52942 89778 53026 90014
rect 53262 89778 88706 90014
rect 88942 89778 89026 90014
rect 89262 89778 124706 90014
rect 124942 89778 125026 90014
rect 125262 89778 160706 90014
rect 160942 89778 161026 90014
rect 161262 89778 196706 90014
rect 196942 89778 197026 90014
rect 197262 89778 232706 90014
rect 232942 89778 233026 90014
rect 233262 89778 268706 90014
rect 268942 89778 269026 90014
rect 269262 89778 304706 90014
rect 304942 89778 305026 90014
rect 305262 89778 340706 90014
rect 340942 89778 341026 90014
rect 341262 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 412706 90014
rect 412942 89778 413026 90014
rect 413262 89778 448706 90014
rect 448942 89778 449026 90014
rect 449262 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 520706 90014
rect 520942 89778 521026 90014
rect 521262 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 592650 90014
rect -8726 89746 592650 89778
rect -8726 86614 592650 86646
rect -8726 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 592650 86294
rect -8726 86026 592650 86058
rect -8726 82894 592650 82926
rect -8726 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 592650 82894
rect -8726 82574 592650 82658
rect -8726 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 592650 82574
rect -8726 82306 592650 82338
rect -8726 79174 592650 79206
rect -8726 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 79426 79174
rect 79662 78938 87867 79174
rect 88103 78938 96308 79174
rect 96544 78938 104749 79174
rect 104985 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 177932 79174
rect 178168 78938 184878 79174
rect 185114 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 191824 79174
rect 192060 78938 198770 79174
rect 199006 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 592650 79174
rect -8726 78854 592650 78938
rect -8726 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 79426 78854
rect 79662 78618 87867 78854
rect 88103 78618 96308 78854
rect 96544 78618 104749 78854
rect 104985 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 177932 78854
rect 178168 78618 184878 78854
rect 185114 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 191824 78854
rect 192060 78618 198770 78854
rect 199006 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 592650 78854
rect -8726 78586 592650 78618
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 75206 75454
rect 75442 75218 83647 75454
rect 83883 75218 92088 75454
rect 92324 75218 100529 75454
rect 100765 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 174459 75454
rect 174695 75218 181405 75454
rect 181641 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 188351 75454
rect 188587 75218 195297 75454
rect 195533 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 75206 75134
rect 75442 74898 83647 75134
rect 83883 74898 92088 75134
rect 92324 74898 100529 75134
rect 100765 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 174459 75134
rect 174695 74898 181405 75134
rect 181641 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 188351 75134
rect 188587 74898 195297 75134
rect 195533 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 65494 592650 65526
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 63866 65494
rect 64102 65258 64186 65494
rect 64422 65258 99866 65494
rect 100102 65258 100186 65494
rect 100422 65258 135866 65494
rect 136102 65258 136186 65494
rect 136422 65258 171866 65494
rect 172102 65258 172186 65494
rect 172422 65258 207866 65494
rect 208102 65258 208186 65494
rect 208422 65258 243866 65494
rect 244102 65258 244186 65494
rect 244422 65258 279866 65494
rect 280102 65258 280186 65494
rect 280422 65258 315866 65494
rect 316102 65258 316186 65494
rect 316422 65258 351866 65494
rect 352102 65258 352186 65494
rect 352422 65258 387866 65494
rect 388102 65258 388186 65494
rect 388422 65258 423866 65494
rect 424102 65258 424186 65494
rect 424422 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect -8726 65174 592650 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 63866 65174
rect 64102 64938 64186 65174
rect 64422 64938 99866 65174
rect 100102 64938 100186 65174
rect 100422 64938 135866 65174
rect 136102 64938 136186 65174
rect 136422 64938 171866 65174
rect 172102 64938 172186 65174
rect 172422 64938 207866 65174
rect 208102 64938 208186 65174
rect 208422 64938 243866 65174
rect 244102 64938 244186 65174
rect 244422 64938 279866 65174
rect 280102 64938 280186 65174
rect 280422 64938 315866 65174
rect 316102 64938 316186 65174
rect 316422 64938 351866 65174
rect 352102 64938 352186 65174
rect 352422 64938 387866 65174
rect 388102 64938 388186 65174
rect 388422 64938 423866 65174
rect 424102 64938 424186 65174
rect 424422 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect -8726 64906 592650 64938
rect -8726 61774 592650 61806
rect -8726 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 24146 61774
rect 24382 61538 24466 61774
rect 24702 61538 60146 61774
rect 60382 61538 60466 61774
rect 60702 61538 96146 61774
rect 96382 61538 96466 61774
rect 96702 61538 132146 61774
rect 132382 61538 132466 61774
rect 132702 61538 168146 61774
rect 168382 61538 168466 61774
rect 168702 61538 204146 61774
rect 204382 61538 204466 61774
rect 204702 61538 240146 61774
rect 240382 61538 240466 61774
rect 240702 61538 276146 61774
rect 276382 61538 276466 61774
rect 276702 61538 312146 61774
rect 312382 61538 312466 61774
rect 312702 61538 348146 61774
rect 348382 61538 348466 61774
rect 348702 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 420146 61774
rect 420382 61538 420466 61774
rect 420702 61538 456146 61774
rect 456382 61538 456466 61774
rect 456702 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 592650 61774
rect -8726 61454 592650 61538
rect -8726 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 24146 61454
rect 24382 61218 24466 61454
rect 24702 61218 60146 61454
rect 60382 61218 60466 61454
rect 60702 61218 96146 61454
rect 96382 61218 96466 61454
rect 96702 61218 132146 61454
rect 132382 61218 132466 61454
rect 132702 61218 168146 61454
rect 168382 61218 168466 61454
rect 168702 61218 204146 61454
rect 204382 61218 204466 61454
rect 204702 61218 240146 61454
rect 240382 61218 240466 61454
rect 240702 61218 276146 61454
rect 276382 61218 276466 61454
rect 276702 61218 312146 61454
rect 312382 61218 312466 61454
rect 312702 61218 348146 61454
rect 348382 61218 348466 61454
rect 348702 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 420146 61454
rect 420382 61218 420466 61454
rect 420702 61218 456146 61454
rect 456382 61218 456466 61454
rect 456702 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 592650 61454
rect -8726 61186 592650 61218
rect -8726 58054 592650 58086
rect -8726 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 56426 58054
rect 56662 57818 56746 58054
rect 56982 57818 92426 58054
rect 92662 57818 92746 58054
rect 92982 57818 128426 58054
rect 128662 57818 128746 58054
rect 128982 57818 164426 58054
rect 164662 57818 164746 58054
rect 164982 57818 200426 58054
rect 200662 57818 200746 58054
rect 200982 57818 236426 58054
rect 236662 57818 236746 58054
rect 236982 57818 272426 58054
rect 272662 57818 272746 58054
rect 272982 57818 308426 58054
rect 308662 57818 308746 58054
rect 308982 57818 344426 58054
rect 344662 57818 344746 58054
rect 344982 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 416426 58054
rect 416662 57818 416746 58054
rect 416982 57818 452426 58054
rect 452662 57818 452746 58054
rect 452982 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 592650 58054
rect -8726 57734 592650 57818
rect -8726 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 56426 57734
rect 56662 57498 56746 57734
rect 56982 57498 92426 57734
rect 92662 57498 92746 57734
rect 92982 57498 128426 57734
rect 128662 57498 128746 57734
rect 128982 57498 164426 57734
rect 164662 57498 164746 57734
rect 164982 57498 200426 57734
rect 200662 57498 200746 57734
rect 200982 57498 236426 57734
rect 236662 57498 236746 57734
rect 236982 57498 272426 57734
rect 272662 57498 272746 57734
rect 272982 57498 308426 57734
rect 308662 57498 308746 57734
rect 308982 57498 344426 57734
rect 344662 57498 344746 57734
rect 344982 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 416426 57734
rect 416662 57498 416746 57734
rect 416982 57498 452426 57734
rect 452662 57498 452746 57734
rect 452982 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 592650 57734
rect -8726 57466 592650 57498
rect -8726 54334 592650 54366
rect -8726 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 52706 54334
rect 52942 54098 53026 54334
rect 53262 54098 88706 54334
rect 88942 54098 89026 54334
rect 89262 54098 124706 54334
rect 124942 54098 125026 54334
rect 125262 54098 160706 54334
rect 160942 54098 161026 54334
rect 161262 54098 196706 54334
rect 196942 54098 197026 54334
rect 197262 54098 232706 54334
rect 232942 54098 233026 54334
rect 233262 54098 268706 54334
rect 268942 54098 269026 54334
rect 269262 54098 304706 54334
rect 304942 54098 305026 54334
rect 305262 54098 340706 54334
rect 340942 54098 341026 54334
rect 341262 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 412706 54334
rect 412942 54098 413026 54334
rect 413262 54098 448706 54334
rect 448942 54098 449026 54334
rect 449262 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 592650 54334
rect -8726 54014 592650 54098
rect -8726 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 52706 54014
rect 52942 53778 53026 54014
rect 53262 53778 88706 54014
rect 88942 53778 89026 54014
rect 89262 53778 124706 54014
rect 124942 53778 125026 54014
rect 125262 53778 160706 54014
rect 160942 53778 161026 54014
rect 161262 53778 196706 54014
rect 196942 53778 197026 54014
rect 197262 53778 232706 54014
rect 232942 53778 233026 54014
rect 233262 53778 268706 54014
rect 268942 53778 269026 54014
rect 269262 53778 304706 54014
rect 304942 53778 305026 54014
rect 305262 53778 340706 54014
rect 340942 53778 341026 54014
rect 341262 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 412706 54014
rect 412942 53778 413026 54014
rect 413262 53778 448706 54014
rect 448942 53778 449026 54014
rect 449262 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 592650 54014
rect -8726 53746 592650 53778
rect -8726 50614 592650 50646
rect -8726 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 592650 50294
rect -8726 50026 592650 50058
rect -8726 46894 592650 46926
rect -8726 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 592650 46894
rect -8726 46574 592650 46658
rect -8726 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 592650 46574
rect -8726 46306 592650 46338
rect -8726 43174 592650 43206
rect -8726 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 592650 43174
rect -8726 42854 592650 42938
rect -8726 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 592650 42854
rect -8726 42586 592650 42618
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 29494 592650 29526
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect -8726 29174 592650 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 592650 25774
rect -8726 25454 592650 25538
rect -8726 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 592650 25454
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 592650 22054
rect -8726 21734 592650 21818
rect -8726 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 592650 21734
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 592650 18334
rect -8726 18014 592650 18098
rect -8726 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 592650 18014
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 592650 14294
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 592650 10894
rect -8726 10574 592650 10658
rect -8726 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 592650 10574
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 592650 7174
rect -8726 6854 592650 6938
rect -8726 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 592650 6854
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use wrapped_channel  wrapped_channel_1
timestamp 0
transform 1 0 70000 0 1 200000
box -10 -52 49800 49828
use wrapped_frequency_counter  wrapped_frequency_counter_2
timestamp 0
transform 1 0 170000 0 1 70000
box -10 -52 29979 49828
use wrapped_rgb_mixer  wrapped_rgb_mixer_3
timestamp 0
transform 1 0 70000 0 1 70000
box -10 -52 35959 41800
use wrapped_simon_game  wrapped_simon_game_4
timestamp 0
transform 1 0 170000 0 1 170000
box -10 -52 59994 59800
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 200068 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 249436 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 177223 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 225473 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 9234 -7654 9854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 -7654 45854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 -7654 81854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 -7654 117854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 -7654 153854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 -7654 189854 92591 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 115001 189854 170068 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 229772 189854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 -7654 225854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 -7654 261854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 -7654 297854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 -7654 333854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 -7654 369854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 -7654 405854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 -7654 441854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 -7654 477854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 -7654 513854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 -7654 549854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 10306 592650 10926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 46306 592650 46926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 82306 592650 82926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 118306 592650 118926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 154306 592650 154926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 190306 592650 190926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 226306 592650 226926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 262306 592650 262926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 298306 592650 298926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 334306 592650 334926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 370306 592650 370926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 406306 592650 406926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 442306 592650 442926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 478306 592650 478926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 514306 592650 514926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 550306 592650 550926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 586306 592650 586926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 622306 592650 622926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 658306 592650 658926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 694306 592650 694926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 16674 -7654 17294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 52674 -7654 53294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 -7654 89294 222319 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 249081 89294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 124674 -7654 125294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 160674 -7654 161294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 -7654 197294 177223 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 225473 197294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 -7654 233294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 -7654 269294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 -7654 305294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 -7654 341294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 376674 -7654 377294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 -7654 413294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 -7654 449294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 -7654 485294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 -7654 521294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 -7654 557294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 17746 592650 18366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 53746 592650 54366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 89746 592650 90366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 125746 592650 126366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 161746 592650 162366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 197746 592650 198366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 233746 592650 234366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 269746 592650 270366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 305746 592650 306366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 341746 592650 342366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 377746 592650 378366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 413746 592650 414366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 449746 592650 450366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 485746 592650 486366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 521746 592650 522366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 557746 592650 558366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 593746 592650 594366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 629746 592650 630366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 665746 592650 666366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 24114 -7654 24734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 60114 -7654 60734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 -7654 96734 70068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 111820 96734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 132114 -7654 132734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 168114 -7654 168734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204114 -7654 204734 177223 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204114 225473 204734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 -7654 240734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 -7654 276734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312114 -7654 312734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 -7654 348734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 384114 -7654 384734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 -7654 420734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 -7654 456734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 -7654 492734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 -7654 528734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 -7654 564734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 25186 592650 25806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 61186 592650 61806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 97186 592650 97806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 133186 592650 133806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 169186 592650 169806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 205186 592650 205806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 241186 592650 241806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 277186 592650 277806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 313186 592650 313806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 349186 592650 349806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 385186 592650 385806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 421186 592650 421806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 457186 592650 457806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 493186 592650 493806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 529186 592650 529806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 565186 592650 565806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 601186 592650 601806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 637186 592650 637806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 673186 592650 673806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 20394 -7654 21014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 56394 -7654 57014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 -7654 93014 70068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 111820 93014 222319 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 249081 93014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 -7654 129014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164394 -7654 165014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 -7654 201014 177223 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 225473 201014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236394 -7654 237014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 -7654 273014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 -7654 309014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 -7654 345014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 380394 -7654 381014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 -7654 417014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 -7654 453014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 -7654 489014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 -7654 525014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 -7654 561014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 21466 592650 22086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 57466 592650 58086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 93466 592650 94086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 129466 592650 130086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 165466 592650 166086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 201466 592650 202086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 237466 592650 238086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 273466 592650 274086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 309466 592650 310086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 345466 592650 346086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 381466 592650 382086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 417466 592650 418086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 453466 592650 454086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 489466 592650 490086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 525466 592650 526086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 561466 592650 562086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 597466 592650 598086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 633466 592650 634086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 669466 592650 670086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 27834 -7654 28454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 -7654 64454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 -7654 100454 70068 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 111820 100454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 -7654 136454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 -7654 172454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 -7654 208454 177223 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 225473 208454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 -7654 244454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 -7654 280454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 315834 -7654 316454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 -7654 352454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 -7654 388454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 -7654 424454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 -7654 460454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 -7654 496454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 -7654 532454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 567834 -7654 568454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 28906 592650 29526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 64906 592650 65526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 100906 592650 101526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 136906 592650 137526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 172906 592650 173526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 208906 592650 209526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 244906 592650 245526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 280906 592650 281526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 316906 592650 317526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 352906 592650 353526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 388906 592650 389526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 424906 592650 425526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 460906 592650 461526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 496906 592650 497526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 532906 592650 533526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 568906 592650 569526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 604906 592650 605526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 640906 592650 641526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 676906 592650 677526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 5514 -7654 6134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 -7654 42134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 -7654 78134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 -7654 114134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 -7654 150134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 -7654 186134 177223 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 225473 186134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 -7654 222134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 -7654 258134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 -7654 294134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 -7654 330134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 -7654 366134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 -7654 402134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 -7654 438134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 -7654 474134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 -7654 510134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 -7654 546134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 581514 -7654 582134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 6586 592650 7206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 42586 592650 43206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 78586 592650 79206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 114586 592650 115206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 150586 592650 151206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 186586 592650 187206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 222586 592650 223206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 258586 592650 259206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 294586 592650 295206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 330586 592650 331206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 366586 592650 367206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 402586 592650 403206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 438586 592650 439206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 474586 592650 475206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 510586 592650 511206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 546586 592650 547206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 582586 592650 583206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 618586 592650 619206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 654586 592650 655206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 690586 592650 691206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 12954 -7654 13574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 -7654 49574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 -7654 85574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 -7654 121574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 -7654 157574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 -7654 193574 177223 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 225473 193574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 -7654 229574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 -7654 265574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 -7654 301574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 -7654 337574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 -7654 373574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 -7654 409574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 -7654 445574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 -7654 481574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 -7654 517574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 -7654 553574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 14026 592650 14646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 50026 592650 50646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 86026 592650 86646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 122026 592650 122646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 158026 592650 158646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 194026 592650 194646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 230026 592650 230646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 266026 592650 266646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 302026 592650 302646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 338026 592650 338646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 374026 592650 374646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 410026 592650 410646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 446026 592650 446646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 482026 592650 482646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 518026 592650 518646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 554026 592650 554646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 590026 592650 590646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 626026 592650 626646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 662026 592650 662646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 698026 592650 698646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
rlabel via4 205088 219336 205088 219336 0 vccd1
rlabel via4 225704 226776 225704 226776 0 vccd2
rlabel via4 89144 90216 89144 90216 0 vdda1
rlabel via4 96584 241656 96584 241656 0 vdda2
rlabel via4 92864 201936 92864 201936 0 vssa1
rlabel via4 208304 173376 208304 173376 0 vssa2
rlabel via4 221984 223056 221984 223056 0 vssd1
rlabel via4 229424 194496 229424 194496 0 vssd2
rlabel metal2 580198 6715 580198 6715 0 io_in[0]
rlabel metal2 97750 250536 97750 250536 0 io_in[10]
rlabel metal2 173190 370532 173190 370532 0 io_in[11]
rlabel metal4 199732 114104 199732 114104 0 io_in[12]
rlabel metal2 93886 199019 93886 199019 0 io_in[13]
rlabel metal2 140806 113849 140806 113849 0 io_in[14]
rlabel metal4 199732 115804 199732 115804 0 io_in[15]
rlabel metal3 231418 174828 231418 174828 0 io_in[16]
rlabel metal2 80086 116382 80086 116382 0 io_in[17]
rlabel metal2 82294 249907 82294 249907 0 io_in[18]
rlabel metal2 299736 703596 299736 703596 0 io_in[19]
rlabel metal2 155894 65382 155894 65382 0 io_in[1]
rlabel metal2 234830 703596 234830 703596 0 io_in[20]
rlabel metal1 67068 218042 67068 218042 0 io_in[21]
rlabel metal2 121486 215883 121486 215883 0 io_in[22]
rlabel metal2 79173 249764 79173 249764 0 io_in[23]
rlabel metal2 76498 250706 76498 250706 0 io_in[24]
rlabel metal2 137310 197880 137310 197880 0 io_in[25]
rlabel metal3 1832 579972 1832 579972 0 io_in[26]
rlabel metal3 1878 527884 1878 527884 0 io_in[27]
rlabel metal3 1556 475660 1556 475660 0 io_in[28]
rlabel metal3 1878 423572 1878 423572 0 io_in[29]
rlabel metal2 233910 76568 233910 76568 0 io_in[2]
rlabel metal3 1970 371348 1970 371348 0 io_in[30]
rlabel metal1 98670 199308 98670 199308 0 io_in[31]
rlabel metal3 1878 267172 1878 267172 0 io_in[32]
rlabel metal3 1832 214948 1832 214948 0 io_in[33]
rlabel metal1 96186 114478 96186 114478 0 io_in[34]
rlabel metal2 113206 250944 113206 250944 0 io_in[35]
rlabel via2 119347 230996 119347 230996 0 io_in[36]
rlabel metal2 114494 251862 114494 251862 0 io_in[37]
rlabel metal2 99038 251590 99038 251590 0 io_in[3]
rlabel metal3 120604 230724 120604 230724 0 io_in[4]
rlabel metal4 199732 118524 199732 118524 0 io_in[5]
rlabel metal2 98670 199512 98670 199512 0 io_in[6]
rlabel metal2 580198 298435 580198 298435 0 io_in[7]
rlabel via2 122498 233291 122498 233291 0 io_in[8]
rlabel metal2 78430 249839 78430 249839 0 io_in[9]
rlabel metal2 96462 185300 96462 185300 0 io_oeb[0]
rlabel metal2 580198 484517 580198 484517 0 io_oeb[10]
rlabel metal4 199732 102884 199732 102884 0 io_oeb[11]
rlabel metal2 121486 214455 121486 214455 0 io_oeb[12]
rlabel metal2 121946 213061 121946 213061 0 io_oeb[13]
rlabel metal3 581908 697204 581908 697204 0 io_oeb[14]
rlabel metal4 119876 249764 119876 249764 0 io_oeb[15]
rlabel metal3 229724 171957 229724 171957 0 io_oeb[16]
rlabel metal2 115874 67048 115874 67048 0 io_oeb[17]
rlabel metal2 213617 229772 213617 229772 0 io_oeb[18]
rlabel metal2 118726 250563 118726 250563 0 io_oeb[19]
rlabel metal2 580198 72369 580198 72369 0 io_oeb[1]
rlabel metal4 199732 97444 199732 97444 0 io_oeb[20]
rlabel metal2 119922 249747 119922 249747 0 io_oeb[21]
rlabel metal2 173926 68690 173926 68690 0 io_oeb[22]
rlabel metal2 94937 249764 94937 249764 0 io_oeb[23]
rlabel metal3 1878 658172 1878 658172 0 io_oeb[24]
rlabel metal2 98762 199546 98762 199546 0 io_oeb[25]
rlabel metal3 230498 216988 230498 216988 0 io_oeb[26]
rlabel metal3 1694 501772 1694 501772 0 io_oeb[27]
rlabel metal3 1740 449548 1740 449548 0 io_oeb[28]
rlabel metal3 120742 232764 120742 232764 0 io_oeb[29]
rlabel metal2 193246 119942 193246 119942 0 io_oeb[2]
rlabel metal3 1832 345372 1832 345372 0 io_oeb[30]
rlabel metal3 1832 293148 1832 293148 0 io_oeb[31]
rlabel metal3 1694 241060 1694 241060 0 io_oeb[32]
rlabel metal3 1878 188836 1878 188836 0 io_oeb[33]
rlabel metal3 1924 136748 1924 136748 0 io_oeb[34]
rlabel metal3 1878 84660 1878 84660 0 io_oeb[35]
rlabel metal3 1556 45492 1556 45492 0 io_oeb[36]
rlabel metal3 1878 6460 1878 6460 0 io_oeb[37]
rlabel metal2 95726 199070 95726 199070 0 io_oeb[3]
rlabel metal2 579738 192185 579738 192185 0 io_oeb[4]
rlabel metal2 580014 231727 580014 231727 0 io_oeb[5]
rlabel metal3 119960 217668 119960 217668 0 io_oeb[6]
rlabel metal2 82938 249890 82938 249890 0 io_oeb[7]
rlabel metal2 173282 68129 173282 68129 0 io_oeb[8]
rlabel metal2 114494 172890 114494 172890 0 io_oeb[9]
rlabel metal1 121670 233206 121670 233206 0 io_out[0]
rlabel via3 120037 95268 120037 95268 0 io_out[10]
rlabel metal3 581954 524484 581954 524484 0 io_out[11]
rlabel metal2 580198 577269 580198 577269 0 io_out[12]
rlabel metal2 140806 174216 140806 174216 0 io_out[13]
rlabel metal3 231587 217940 231587 217940 0 io_out[14]
rlabel metal2 542386 479883 542386 479883 0 io_out[15]
rlabel metal2 120106 94860 120106 94860 0 io_out[16]
rlabel metal2 116426 250519 116426 250519 0 io_out[17]
rlabel metal2 347806 435377 347806 435377 0 io_out[18]
rlabel metal3 170292 198409 170292 198409 0 io_out[19]
rlabel metal2 120014 250784 120014 250784 0 io_out[1]
rlabel metal2 137402 116960 137402 116960 0 io_out[20]
rlabel metal2 153870 236878 153870 236878 0 io_out[21]
rlabel metal2 133814 65858 133814 65858 0 io_out[22]
rlabel metal1 24932 699686 24932 699686 0 io_out[23]
rlabel metal3 1924 671228 1924 671228 0 io_out[24]
rlabel metal3 1740 619140 1740 619140 0 io_out[25]
rlabel metal3 1878 566916 1878 566916 0 io_out[26]
rlabel metal2 134642 115634 134642 115634 0 io_out[27]
rlabel metal3 1786 462604 1786 462604 0 io_out[28]
rlabel metal3 1878 410516 1878 410516 0 io_out[29]
rlabel metal2 580198 99433 580198 99433 0 io_out[2]
rlabel metal3 1924 358428 1924 358428 0 io_out[30]
rlabel metal2 3772 229080 3772 229080 0 io_out[31]
rlabel metal3 1740 254116 1740 254116 0 io_out[32]
rlabel metal3 230912 178228 230912 178228 0 io_out[33]
rlabel metal3 229900 219028 229900 219028 0 io_out[34]
rlabel metal3 1970 97580 1970 97580 0 io_out[35]
rlabel metal3 1924 58548 1924 58548 0 io_out[36]
rlabel metal3 1924 19380 1924 19380 0 io_out[37]
rlabel metal3 581908 139332 581908 139332 0 io_out[3]
rlabel metal3 120604 229228 120604 229228 0 io_out[4]
rlabel metal2 178434 120843 178434 120843 0 io_out[5]
rlabel metal2 118358 250536 118358 250536 0 io_out[6]
rlabel metal2 580198 311967 580198 311967 0 io_out[7]
rlabel metal2 579830 364735 579830 364735 0 io_out[8]
rlabel metal2 580198 418217 580198 418217 0 io_out[9]
rlabel metal2 129161 340 129161 340 0 la_data_in[1]
rlabel metal2 132756 16560 132756 16560 0 la_data_in[2]
rlabel metal3 230820 179588 230820 179588 0 la_data_in[32]
rlabel metal2 89930 198900 89930 198900 0 la_data_in[33]
rlabel metal2 179078 69642 179078 69642 0 la_data_in[34]
rlabel metal1 159068 111826 159068 111826 0 la_data_in[35]
rlabel metal2 193890 120894 193890 120894 0 la_data_in[36]
rlabel metal4 199732 99756 199732 99756 0 la_data_in[37]
rlabel metal2 193699 229772 193699 229772 0 la_data_in[38]
rlabel metal2 157366 198832 157366 198832 0 la_data_in[39]
rlabel metal2 136482 1894 136482 1894 0 la_data_in[3]
rlabel metal2 194987 229772 194987 229772 0 la_data_in[40]
rlabel metal2 271025 340 271025 340 0 la_data_in[41]
rlabel metal2 274850 2676 274850 2676 0 la_data_in[42]
rlabel metal2 118174 78710 118174 78710 0 la_data_in[43]
rlabel metal1 154928 115634 154928 115634 0 la_data_in[44]
rlabel metal2 196873 70244 196873 70244 0 la_data_in[45]
rlabel metal2 288742 16560 288742 16560 0 la_data_in[46]
rlabel metal2 158102 180064 158102 180064 0 la_data_in[47]
rlabel metal2 101614 250740 101614 250740 0 la_data_in[48]
rlabel metal2 93886 251420 93886 251420 0 la_data_in[49]
rlabel metal2 139833 340 139833 340 0 la_data_in[4]
rlabel metal2 113574 69275 113574 69275 0 la_data_in[50]
rlabel metal2 191169 229772 191169 229772 0 la_data_in[51]
rlabel metal2 310033 340 310033 340 0 la_data_in[52]
rlabel metal2 119002 250502 119002 250502 0 la_data_in[53]
rlabel metal1 116978 121482 116978 121482 0 la_data_in[54]
rlabel metal2 168130 64328 168130 64328 0 la_data_in[55]
rlabel metal2 156722 168742 156722 168742 0 la_data_in[56]
rlabel metal2 327566 16560 327566 16560 0 la_data_in[57]
rlabel metal3 230912 173468 230912 173468 0 la_data_in[58]
rlabel metal2 98946 199206 98946 199206 0 la_data_in[59]
rlabel metal2 64262 105672 64262 105672 0 la_data_in[60]
rlabel metal2 171251 229772 171251 229772 0 la_data_in[61]
rlabel metal2 345545 340 345545 340 0 la_data_in[62]
rlabel metal3 199364 69889 199364 69889 0 la_data_in[63]
rlabel metal2 176219 70244 176219 70244 0 la_data_out[32]
rlabel metal1 67436 114274 67436 114274 0 la_data_out[33]
rlabel metal2 90666 191386 90666 191386 0 la_data_out[34]
rlabel metal2 251206 1911 251206 1911 0 la_data_out[35]
rlabel metal2 254465 340 254465 340 0 la_data_out[36]
rlabel metal2 173190 39655 173190 39655 0 la_data_out[37]
rlabel metal4 199732 96764 199732 96764 0 la_data_out[38]
rlabel metal2 265374 1758 265374 1758 0 la_data_out[39]
rlabel metal1 118818 194922 118818 194922 0 la_data_out[40]
rlabel metal2 117070 250604 117070 250604 0 la_data_out[41]
rlabel metal1 117254 82824 117254 82824 0 la_data_out[42]
rlabel metal2 94622 183294 94622 183294 0 la_data_out[43]
rlabel metal4 199732 117164 199732 117164 0 la_data_out[44]
rlabel metal2 74566 250638 74566 250638 0 la_data_out[45]
rlabel metal2 97106 250706 97106 250706 0 la_data_out[46]
rlabel metal2 293473 340 293473 340 0 la_data_out[47]
rlabel metal2 122038 214829 122038 214829 0 la_data_out[48]
rlabel metal1 119278 193698 119278 193698 0 la_data_out[49]
rlabel metal2 75854 251532 75854 251532 0 la_data_out[50]
rlabel metal1 121854 212466 121854 212466 0 la_data_out[51]
rlabel metal2 311466 1911 311466 1911 0 la_data_out[52]
rlabel metal4 199732 115124 199732 115124 0 la_data_out[53]
rlabel metal2 100326 250502 100326 250502 0 la_data_out[54]
rlabel metal2 116702 183872 116702 183872 0 la_data_out[55]
rlabel metal3 119508 218741 119508 218741 0 la_data_out[56]
rlabel metal2 328985 340 328985 340 0 la_data_out[57]
rlabel metal3 230866 176188 230866 176188 0 la_data_out[58]
rlabel metal2 117990 250478 117990 250478 0 la_data_out[59]
rlabel metal2 115322 176528 115322 176528 0 la_data_out[60]
rlabel metal2 174570 37512 174570 37512 0 la_data_out[61]
rlabel metal3 120742 213044 120742 213044 0 la_data_out[62]
rlabel metal3 121064 248948 121064 248948 0 la_data_out[63]
rlabel metal2 118174 75650 118174 75650 0 la_oenb[32]
rlabel metal2 177291 70244 177291 70244 0 la_oenb[33]
rlabel metal2 248623 340 248623 340 0 la_oenb[34]
rlabel metal2 118818 250818 118818 250818 0 la_oenb[35]
rlabel metal2 155250 122366 155250 122366 0 la_oenb[36]
rlabel metal2 120934 241468 120934 241468 0 la_oenb[37]
rlabel metal2 77786 251896 77786 251896 0 la_oenb[38]
rlabel metal2 197754 69506 197754 69506 0 la_oenb[39]
rlabel metal2 269606 16560 269606 16560 0 la_oenb[40]
rlabel metal2 273463 340 273463 340 0 la_oenb[41]
rlabel metal2 119186 249016 119186 249016 0 la_oenb[42]
rlabel metal1 68632 233886 68632 233886 0 la_oenb[43]
rlabel metal2 64722 104890 64722 104890 0 la_oenb[44]
rlabel metal2 287585 340 287585 340 0 la_oenb[45]
rlabel metal2 291318 16560 291318 16560 0 la_oenb[46]
rlabel metal2 113298 132090 113298 132090 0 la_oenb[47]
rlabel metal1 66838 97954 66838 97954 0 la_oenb[48]
rlabel metal2 175214 230510 175214 230510 0 la_oenb[49]
rlabel metal2 177790 120282 177790 120282 0 la_oenb[50]
rlabel metal2 309074 1860 309074 1860 0 la_oenb[51]
rlabel metal2 312662 1996 312662 1996 0 la_oenb[52]
rlabel metal2 102258 250876 102258 250876 0 la_oenb[53]
rlabel metal2 177146 120588 177146 120588 0 la_oenb[54]
rlabel metal2 94438 197642 94438 197642 0 la_oenb[55]
rlabel metal1 98532 115906 98532 115906 0 la_oenb[56]
rlabel metal3 121087 210188 121087 210188 0 la_oenb[57]
rlabel metal2 119186 251277 119186 251277 0 la_oenb[58]
rlabel metal2 122314 235025 122314 235025 0 la_oenb[59]
rlabel metal2 61870 133450 61870 133450 0 la_oenb[60]
rlabel metal2 115874 68272 115874 68272 0 la_oenb[61]
rlabel via2 122498 234651 122498 234651 0 la_oenb[62]
rlabel metal2 98302 197676 98302 197676 0 la_oenb[63]
rlabel metal2 598 1588 598 1588 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
